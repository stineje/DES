module exp_d(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b100000;
				6'b000001 : out = 8'b000001;
				6'b000010 : out = 8'b000010;
				6'b000011 : out = 8'b000011;
				6'b000100 : out = 8'b000100;
				6'b000101 : out = 8'b000101;
				6'b000110 : out = 8'b000100;
				6'b000111 : out = 8'b000101;
				6'b001000 : out = 8'b000110;
				6'b001001 : out = 8'b000111;
				6'b001010 : out = 8'b001000;
				6'b001011 : out = 8'b001001;
				6'b001100 : out = 8'b001000;
				6'b001101 : out = 8'b001001;
				6'b001110 : out = 8'b001010;
				6'b001111 : out = 8'b001011;
				6'b010000 : out = 8'b001100;
				6'b010001 : out = 8'b001101;
				6'b010010 : out = 8'b001100;
				6'b010011 : out = 8'b001101;
				6'b010100 : out = 8'b001110;
				6'b010101 : out = 8'b001111;
				6'b010110 : out = 8'b010000;
				6'b010111 : out = 8'b010001;
				6'b011000 : out = 8'b010000;
				6'b011001 : out = 8'b010001;
				6'b011010 : out = 8'b010010;
				6'b011011 : out = 8'b010011;
				6'b011100 : out = 8'b010100;
				6'b011101 : out = 8'b010101;
				6'b011110 : out = 8'b010100;
				6'b011111 : out = 8'b010101;
				6'b100000 : out = 8'b010110;
				6'b100001 : out = 8'b010111;
				6'b100010 : out = 8'b011000;
				6'b100011 : out = 8'b011001;
				6'b100100 : out = 8'b011000;
				6'b100101 : out = 8'b011001;
				6'b100110 : out = 8'b011010;
				6'b100111 : out = 8'b011011;
				6'b101000 : out = 8'b011100;
				6'b101001 : out = 8'b011101;
				6'b101010 : out = 8'b011100;
				6'b101011 : out = 8'b011101;
				6'b101100 : out = 8'b011110;
				6'b101101 : out = 8'b011111;
				6'b101110 : out = 8'b100000;
				6'b101111 : out = 8'b000001;
			endcase
		  end

endmodule

module final_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0101000;
				7'b0000001 : out = 8'b0001000;
				7'b0000010 : out = 8'b0110000;
				7'b0000011 : out = 8'b0010000;
				7'b0000100 : out = 8'b0111000;
				7'b0000101 : out = 8'b0011000;
				7'b0000110 : out = 8'b1000000;
				7'b0000111 : out = 8'b0100000;
				7'b0001000 : out = 8'b0100111;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0101111;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0110111;
				7'b0001101 : out = 8'b0010111;
				7'b0001110 : out = 8'b0111111;
				7'b0001111 : out = 8'b0011111;
				7'b0010000 : out = 8'b0100110;
				7'b0010001 : out = 8'b0000110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0001110;
				7'b0010100 : out = 8'b0110110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0111110;
				7'b0010111 : out = 8'b0011110;
				7'b0011000 : out = 8'b0100101;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0101101;
				7'b0011011 : out = 8'b0001101;
				7'b0011100 : out = 8'b0110101;
				7'b0011101 : out = 8'b0010101;
				7'b0011110 : out = 8'b0111101;
				7'b0011111 : out = 8'b0011101;
				7'b0100000 : out = 8'b0100100;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0101100;
				7'b0100011 : out = 8'b0001100;
				7'b0100100 : out = 8'b0110100;
				7'b0100101 : out = 8'b0010100;
				7'b0100110 : out = 8'b0111100;
				7'b0100111 : out = 8'b0011100;
				7'b0101000 : out = 8'b0100011;
				7'b0101001 : out = 8'b0000011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0001011;
				7'b0101100 : out = 8'b0110011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0111011;
				7'b0101111 : out = 8'b0011011;
				7'b0110000 : out = 8'b0100010;
				7'b0110001 : out = 8'b0000010;
				7'b0110010 : out = 8'b0101010;
				7'b0110011 : out = 8'b0001010;
				7'b0110100 : out = 8'b0110010;
				7'b0110101 : out = 8'b0010010;
				7'b0110110 : out = 8'b0111010;
				7'b0110111 : out = 8'b0011010;
				7'b0111000 : out = 8'b0100001;
				7'b0111001 : out = 8'b0000001;
				7'b0111010 : out = 8'b0101001;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0110001;
				7'b0111101 : out = 8'b0010001;
				7'b0111110 : out = 8'b0111001;
				7'b0111111 : out = 8'b0011001;
			endcase
		  end

endmodule

module initial_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0111010;
				7'b0000001 : out = 8'b0110010;
				7'b0000010 : out = 8'b0101010;
				7'b0000011 : out = 8'b0100010;
				7'b0000100 : out = 8'b0011010;
				7'b0000101 : out = 8'b0010010;
				7'b0000110 : out = 8'b0001010;
				7'b0000111 : out = 8'b0000010;
				7'b0001000 : out = 8'b0111100;
				7'b0001001 : out = 8'b0110100;
				7'b0001010 : out = 8'b0101100;
				7'b0001011 : out = 8'b0100100;
				7'b0001100 : out = 8'b0011100;
				7'b0001101 : out = 8'b0010100;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000100;
				7'b0010000 : out = 8'b0111110;
				7'b0010001 : out = 8'b0110110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0100110;
				7'b0010100 : out = 8'b0011110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0001110;
				7'b0010111 : out = 8'b0000110;
				7'b0011000 : out = 8'b1000000;
				7'b0011001 : out = 8'b0111000;
				7'b0011010 : out = 8'b0110000;
				7'b0011011 : out = 8'b0101000;
				7'b0011100 : out = 8'b0100000;
				7'b0011101 : out = 8'b0011000;
				7'b0011110 : out = 8'b0010000;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0111001;
				7'b0100001 : out = 8'b0110001;
				7'b0100010 : out = 8'b0101001;
				7'b0100011 : out = 8'b0100001;
				7'b0100100 : out = 8'b0011001;
				7'b0100101 : out = 8'b0010001;
				7'b0100110 : out = 8'b0001001;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0111011;
				7'b0101001 : out = 8'b0110011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0100011;
				7'b0101100 : out = 8'b0011011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000011;
				7'b0110000 : out = 8'b0111101;
				7'b0110001 : out = 8'b0110101;
				7'b0110010 : out = 8'b0101101;
				7'b0110011 : out = 8'b0100101;
				7'b0110100 : out = 8'b0011101;
				7'b0110101 : out = 8'b0010101;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0000101;
				7'b0111000 : out = 8'b0111111;
				7'b0111001 : out = 8'b0110111;
				7'b0111010 : out = 8'b0101111;
				7'b0111011 : out = 8'b0100111;
				7'b0111100 : out = 8'b0011111;
				7'b0111101 : out = 8'b0010111;
				7'b0111110 : out = 8'b0001111;
				7'b0111111 : out = 8'b0000111;
			endcase
		  end

endmodule

module per(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b010000;
				6'b000001 : out = 8'b000111;
				6'b000010 : out = 8'b010100;
				6'b000011 : out = 8'b010101;
				6'b000100 : out = 8'b011101;
				6'b000101 : out = 8'b001100;
				6'b000110 : out = 8'b011100;
				6'b000111 : out = 8'b010001;
				6'b001000 : out = 8'b000001;
				6'b001001 : out = 8'b001111;
				6'b001010 : out = 8'b010111;
				6'b001011 : out = 8'b011010;
				6'b001100 : out = 8'b000101;
				6'b001101 : out = 8'b010010;
				6'b001110 : out = 8'b011111;
				6'b001111 : out = 8'b001010;
				6'b010000 : out = 8'b000010;
				6'b010001 : out = 8'b001000;
				6'b010010 : out = 8'b011000;
				6'b010011 : out = 8'b001110;
				6'b010100 : out = 8'b100000;
				6'b010101 : out = 8'b011011;
				6'b010110 : out = 8'b000011;
				6'b010111 : out = 8'b001001;
				6'b011000 : out = 8'b010011;
				6'b011001 : out = 8'b001101;
				6'b011010 : out = 8'b011110;
				6'b011011 : out = 8'b000110;
				6'b011100 : out = 8'b010110;
				6'b011101 : out = 8'b001011;
				6'b011110 : out = 8'b000100;
				6'b011111 : out = 8'b011001;
			endcase
		  end

endmodule

module sbox_0(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001110;
				7'b0000001 : out = 8'b0000100;
				7'b0000010 : out = 8'b0001101;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000010;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001010;
				7'b0001010 : out = 8'b0000110;
				7'b0001011 : out = 8'b0001100;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001001;
				7'b0001110 : out = 8'b0000000;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000000;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000111;
				7'b0010011 : out = 8'b0000100;
				7'b0010100 : out = 8'b0001110;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0001010;
				7'b0011001 : out = 8'b0000110;
				7'b0011010 : out = 8'b0001100;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0001001;
				7'b0011101 : out = 8'b0000101;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000001;
				7'b0100010 : out = 8'b0001110;
				7'b0100011 : out = 8'b0001000;
				7'b0100100 : out = 8'b0001101;
				7'b0100101 : out = 8'b0000110;
				7'b0100110 : out = 8'b0000010;
				7'b0100111 : out = 8'b0001011;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001100;
				7'b0101010 : out = 8'b0001001;
				7'b0101011 : out = 8'b0000111;
				7'b0101100 : out = 8'b0000011;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0000000;
				7'b0110000 : out = 8'b0001111;
				7'b0110001 : out = 8'b0001100;
				7'b0110010 : out = 8'b0001000;
				7'b0110011 : out = 8'b0000010;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0000001;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000101;
				7'b0111001 : out = 8'b0001011;
				7'b0111010 : out = 8'b0000011;
				7'b0111011 : out = 8'b0001110;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule

module sbox_1(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001111;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001011;
				7'b0000110 : out = 8'b0000011;
				7'b0000111 : out = 8'b0000100;
				7'b0001000 : out = 8'b0001001;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0000010;
				7'b0001011 : out = 8'b0001101;
				7'b0001100 : out = 8'b0001100;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001010;
				7'b0010000 : out = 8'b0000011;
				7'b0010001 : out = 8'b0001101;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0001111;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001000;
				7'b0010111 : out = 8'b0001110;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0000001;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000110;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001011;
				7'b0011111 : out = 8'b0000101;
				7'b0100000 : out = 8'b0000000;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0000111;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0000100;
				7'b0100110 : out = 8'b0001101;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0000101;
				7'b0101001 : out = 8'b0001000;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000110;
				7'b0101100 : out = 8'b0001001;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000010;
				7'b0101111 : out = 8'b0001111;
				7'b0110000 : out = 8'b0001101;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001010;
				7'b0110011 : out = 8'b0000001;
				7'b0110100 : out = 8'b0000011;
				7'b0110101 : out = 8'b0001111;
				7'b0110110 : out = 8'b0000100;
				7'b0110111 : out = 8'b0000010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0000110;
				7'b0111010 : out = 8'b0000111;
				7'b0111011 : out = 8'b0001100;
				7'b0111100 : out = 8'b0000000;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0001110;
				7'b0111111 : out = 8'b0001001;
			endcase
		  end

endmodule

module sbox_2(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001010;
				7'b0000001 : out = 8'b0000000;
				7'b0000010 : out = 8'b0001001;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0000011;
				7'b0000110 : out = 8'b0001111;
				7'b0000111 : out = 8'b0000101;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0001100;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0000100;
				7'b0001110 : out = 8'b0000010;
				7'b0001111 : out = 8'b0001000;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000111;
				7'b0010010 : out = 8'b0000000;
				7'b0010011 : out = 8'b0001001;
				7'b0010100 : out = 8'b0000011;
				7'b0010101 : out = 8'b0000100;
				7'b0010110 : out = 8'b0000110;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0000010;
				7'b0011001 : out = 8'b0001000;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0001100;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0001111;
				7'b0011111 : out = 8'b0000001;
				7'b0100000 : out = 8'b0001101;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0001001;
				7'b0100100 : out = 8'b0001000;
				7'b0100101 : out = 8'b0001111;
				7'b0100110 : out = 8'b0000011;
				7'b0100111 : out = 8'b0000000;
				7'b0101000 : out = 8'b0001011;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000010;
				7'b0101011 : out = 8'b0001100;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0001110;
				7'b0101111 : out = 8'b0000111;
				7'b0110000 : out = 8'b0000001;
				7'b0110001 : out = 8'b0001010;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0000000;
				7'b0110100 : out = 8'b0000110;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000100;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0001110;
				7'b0111011 : out = 8'b0000011;
				7'b0111100 : out = 8'b0001011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule

module sbox_3(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000111;
				7'b0000001 : out = 8'b0001101;
				7'b0000010 : out = 8'b0001110;
				7'b0000011 : out = 8'b0000011;
				7'b0000100 : out = 8'b0000000;
				7'b0000101 : out = 8'b0000110;
				7'b0000110 : out = 8'b0001001;
				7'b0000111 : out = 8'b0001010;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0000010;
				7'b0001010 : out = 8'b0001000;
				7'b0001011 : out = 8'b0000101;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0001100;
				7'b0001110 : out = 8'b0000100;
				7'b0001111 : out = 8'b0001111;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0001000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000101;
				7'b0010100 : out = 8'b0000110;
				7'b0010101 : out = 8'b0001111;
				7'b0010110 : out = 8'b0000000;
				7'b0010111 : out = 8'b0000011;
				7'b0011000 : out = 8'b0000100;
				7'b0011001 : out = 8'b0000111;
				7'b0011010 : out = 8'b0000010;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000001;
				7'b0011101 : out = 8'b0001010;
				7'b0011110 : out = 8'b0001110;
				7'b0011111 : out = 8'b0001001;
				7'b0100000 : out = 8'b0001010;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0001001;
				7'b0100011 : out = 8'b0000000;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0001011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001101;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000011;
				7'b0101011 : out = 8'b0001110;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0000010;
				7'b0101110 : out = 8'b0001000;
				7'b0101111 : out = 8'b0000100;
				7'b0110000 : out = 8'b0000011;
				7'b0110001 : out = 8'b0001111;
				7'b0110010 : out = 8'b0000000;
				7'b0110011 : out = 8'b0000110;
				7'b0110100 : out = 8'b0001010;
				7'b0110101 : out = 8'b0000001;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0001000;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000100;
				7'b0111010 : out = 8'b0000101;
				7'b0111011 : out = 8'b0001011;
				7'b0111100 : out = 8'b0001100;
				7'b0111101 : out = 8'b0000111;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001110;
			endcase
		  end

endmodule

module sbox_4(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000010;
				7'b0000001 : out = 8'b0001100;
				7'b0000010 : out = 8'b0000100;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000111;
				7'b0000101 : out = 8'b0001010;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000110;
				7'b0001000 : out = 8'b0001000;
				7'b0001001 : out = 8'b0000101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0001101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001110;
				7'b0001111 : out = 8'b0001001;
				7'b0010000 : out = 8'b0001110;
				7'b0010001 : out = 8'b0001011;
				7'b0010010 : out = 8'b0000010;
				7'b0010011 : out = 8'b0001100;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0000111;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0000101;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0001111;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000011;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000010;
				7'b0100010 : out = 8'b0000001;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0001101;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001000;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001001;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000101;
				7'b0101100 : out = 8'b0000110;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000000;
				7'b0101111 : out = 8'b0001110;
				7'b0110000 : out = 8'b0001011;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001100;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0001110;
				7'b0110110 : out = 8'b0000010;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0000110;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000100;
				7'b0111110 : out = 8'b0000101;
				7'b0111111 : out = 8'b0000011;
			endcase
		  end

endmodule

module sbox_5(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001100;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001010;
				7'b0000011 : out = 8'b0001111;
				7'b0000100 : out = 8'b0001001;
				7'b0000101 : out = 8'b0000010;
				7'b0000110 : out = 8'b0000110;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000000;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0000100;
				7'b0001100 : out = 8'b0001110;
				7'b0001101 : out = 8'b0000111;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001011;
				7'b0010000 : out = 8'b0001010;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000010;
				7'b0010100 : out = 8'b0000111;
				7'b0010101 : out = 8'b0001100;
				7'b0010110 : out = 8'b0001001;
				7'b0010111 : out = 8'b0000101;
				7'b0011000 : out = 8'b0000110;
				7'b0011001 : out = 8'b0000001;
				7'b0011010 : out = 8'b0001101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0001001;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0001111;
				7'b0100011 : out = 8'b0000101;
				7'b0100100 : out = 8'b0000010;
				7'b0100101 : out = 8'b0001000;
				7'b0100110 : out = 8'b0001100;
				7'b0100111 : out = 8'b0000011;
				7'b0101000 : out = 8'b0000111;
				7'b0101001 : out = 8'b0000000;
				7'b0101010 : out = 8'b0000100;
				7'b0101011 : out = 8'b0001010;
				7'b0101100 : out = 8'b0000001;
				7'b0101101 : out = 8'b0001101;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000110;
				7'b0110000 : out = 8'b0000100;
				7'b0110001 : out = 8'b0000011;
				7'b0110010 : out = 8'b0000010;
				7'b0110011 : out = 8'b0001100;
				7'b0110100 : out = 8'b0001001;
				7'b0110101 : out = 8'b0000101;
				7'b0110110 : out = 8'b0001111;
				7'b0110111 : out = 8'b0001010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0001110;
				7'b0111010 : out = 8'b0000001;
				7'b0111011 : out = 8'b0000111;
				7'b0111100 : out = 8'b0000110;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0001000;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule

module sbox_6(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000100;
				7'b0000001 : out = 8'b0001011;
				7'b0000010 : out = 8'b0000010;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0001111;
				7'b0000101 : out = 8'b0000000;
				7'b0000110 : out = 8'b0001000;
				7'b0000111 : out = 8'b0001101;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001100;
				7'b0001010 : out = 8'b0001001;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001010;
				7'b0001110 : out = 8'b0000110;
				7'b0001111 : out = 8'b0000001;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0001001;
				7'b0010110 : out = 8'b0000001;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0001110;
				7'b0011001 : out = 8'b0000011;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000010;
				7'b0011101 : out = 8'b0001111;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000001;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0001011;
				7'b0100011 : out = 8'b0001101;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0000011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001110;
				7'b0101000 : out = 8'b0001010;
				7'b0101001 : out = 8'b0001111;
				7'b0101010 : out = 8'b0000110;
				7'b0101011 : out = 8'b0001000;
				7'b0101100 : out = 8'b0000000;
				7'b0101101 : out = 8'b0000101;
				7'b0101110 : out = 8'b0001001;
				7'b0101111 : out = 8'b0000010;
				7'b0110000 : out = 8'b0000110;
				7'b0110001 : out = 8'b0001011;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0001000;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0000100;
				7'b0110110 : out = 8'b0001010;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000101;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001111;
				7'b0111100 : out = 8'b0001110;
				7'b0111101 : out = 8'b0000010;
				7'b0111110 : out = 8'b0000011;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule

module sbox_7(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001101;
				7'b0000001 : out = 8'b0000010;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0000100;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000001;
				7'b0001000 : out = 8'b0001010;
				7'b0001001 : out = 8'b0001001;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001110;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000001;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0001101;
				7'b0010011 : out = 8'b0001000;
				7'b0010100 : out = 8'b0001010;
				7'b0010101 : out = 8'b0000011;
				7'b0010110 : out = 8'b0000111;
				7'b0010111 : out = 8'b0000100;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0000110;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001110;
				7'b0011110 : out = 8'b0001001;
				7'b0011111 : out = 8'b0000010;
				7'b0100000 : out = 8'b0000111;
				7'b0100001 : out = 8'b0001011;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0000001;
				7'b0100100 : out = 8'b0001001;
				7'b0100101 : out = 8'b0001100;
				7'b0100110 : out = 8'b0001110;
				7'b0100111 : out = 8'b0000010;
				7'b0101000 : out = 8'b0000000;
				7'b0101001 : out = 8'b0000110;
				7'b0101010 : out = 8'b0001010;
				7'b0101011 : out = 8'b0001101;
				7'b0101100 : out = 8'b0001111;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0001000;
				7'b0110000 : out = 8'b0000010;
				7'b0110001 : out = 8'b0000001;
				7'b0110010 : out = 8'b0001110;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001010;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0001111;
				7'b0111001 : out = 8'b0001100;
				7'b0111010 : out = 8'b0001001;
				7'b0111011 : out = 8'b0000000;
				7'b0111100 : out = 8'b0000011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001011;
			endcase
		  end

endmodule

module exp_d(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b100000;
				6'b000001 : out = 8'b000001;
				6'b000010 : out = 8'b000010;
				6'b000011 : out = 8'b000011;
				6'b000100 : out = 8'b000100;
				6'b000101 : out = 8'b000101;
				6'b000110 : out = 8'b000100;
				6'b000111 : out = 8'b000101;
				6'b001000 : out = 8'b000110;
				6'b001001 : out = 8'b000111;
				6'b001010 : out = 8'b001000;
				6'b001011 : out = 8'b001001;
				6'b001100 : out = 8'b001000;
				6'b001101 : out = 8'b001001;
				6'b001110 : out = 8'b001010;
				6'b001111 : out = 8'b001011;
				6'b010000 : out = 8'b001100;
				6'b010001 : out = 8'b001101;
				6'b010010 : out = 8'b001100;
				6'b010011 : out = 8'b001101;
				6'b010100 : out = 8'b001110;
				6'b010101 : out = 8'b001111;
				6'b010110 : out = 8'b010000;
				6'b010111 : out = 8'b010001;
				6'b011000 : out = 8'b010000;
				6'b011001 : out = 8'b010001;
				6'b011010 : out = 8'b010010;
				6'b011011 : out = 8'b010011;
				6'b011100 : out = 8'b010100;
				6'b011101 : out = 8'b010101;
				6'b011110 : out = 8'b010100;
				6'b011111 : out = 8'b010101;
				6'b100000 : out = 8'b010110;
				6'b100001 : out = 8'b010111;
				6'b100010 : out = 8'b011000;
				6'b100011 : out = 8'b011001;
				6'b100100 : out = 8'b011000;
				6'b100101 : out = 8'b011001;
				6'b100110 : out = 8'b011010;
				6'b100111 : out = 8'b011011;
				6'b101000 : out = 8'b011100;
				6'b101001 : out = 8'b011101;
				6'b101010 : out = 8'b011100;
				6'b101011 : out = 8'b011101;
				6'b101100 : out = 8'b011110;
				6'b101101 : out = 8'b011111;
				6'b101110 : out = 8'b100000;
				6'b101111 : out = 8'b000001;
			endcase
		  end

endmodule

module final_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0101000;
				7'b0000001 : out = 8'b0001000;
				7'b0000010 : out = 8'b0110000;
				7'b0000011 : out = 8'b0010000;
				7'b0000100 : out = 8'b0111000;
				7'b0000101 : out = 8'b0011000;
				7'b0000110 : out = 8'b1000000;
				7'b0000111 : out = 8'b0100000;
				7'b0001000 : out = 8'b0100111;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0101111;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0110111;
				7'b0001101 : out = 8'b0010111;
				7'b0001110 : out = 8'b0111111;
				7'b0001111 : out = 8'b0011111;
				7'b0010000 : out = 8'b0100110;
				7'b0010001 : out = 8'b0000110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0001110;
				7'b0010100 : out = 8'b0110110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0111110;
				7'b0010111 : out = 8'b0011110;
				7'b0011000 : out = 8'b0100101;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0101101;
				7'b0011011 : out = 8'b0001101;
				7'b0011100 : out = 8'b0110101;
				7'b0011101 : out = 8'b0010101;
				7'b0011110 : out = 8'b0111101;
				7'b0011111 : out = 8'b0011101;
				7'b0100000 : out = 8'b0100100;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0101100;
				7'b0100011 : out = 8'b0001100;
				7'b0100100 : out = 8'b0110100;
				7'b0100101 : out = 8'b0010100;
				7'b0100110 : out = 8'b0111100;
				7'b0100111 : out = 8'b0011100;
				7'b0101000 : out = 8'b0100011;
				7'b0101001 : out = 8'b0000011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0001011;
				7'b0101100 : out = 8'b0110011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0111011;
				7'b0101111 : out = 8'b0011011;
				7'b0110000 : out = 8'b0100010;
				7'b0110001 : out = 8'b0000010;
				7'b0110010 : out = 8'b0101010;
				7'b0110011 : out = 8'b0001010;
				7'b0110100 : out = 8'b0110010;
				7'b0110101 : out = 8'b0010010;
				7'b0110110 : out = 8'b0111010;
				7'b0110111 : out = 8'b0011010;
				7'b0111000 : out = 8'b0100001;
				7'b0111001 : out = 8'b0000001;
				7'b0111010 : out = 8'b0101001;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0110001;
				7'b0111101 : out = 8'b0010001;
				7'b0111110 : out = 8'b0111001;
				7'b0111111 : out = 8'b0011001;
			endcase
		  end

endmodule

module initial_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0111010;
				7'b0000001 : out = 8'b0110010;
				7'b0000010 : out = 8'b0101010;
				7'b0000011 : out = 8'b0100010;
				7'b0000100 : out = 8'b0011010;
				7'b0000101 : out = 8'b0010010;
				7'b0000110 : out = 8'b0001010;
				7'b0000111 : out = 8'b0000010;
				7'b0001000 : out = 8'b0111100;
				7'b0001001 : out = 8'b0110100;
				7'b0001010 : out = 8'b0101100;
				7'b0001011 : out = 8'b0100100;
				7'b0001100 : out = 8'b0011100;
				7'b0001101 : out = 8'b0010100;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000100;
				7'b0010000 : out = 8'b0111110;
				7'b0010001 : out = 8'b0110110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0100110;
				7'b0010100 : out = 8'b0011110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0001110;
				7'b0010111 : out = 8'b0000110;
				7'b0011000 : out = 8'b1000000;
				7'b0011001 : out = 8'b0111000;
				7'b0011010 : out = 8'b0110000;
				7'b0011011 : out = 8'b0101000;
				7'b0011100 : out = 8'b0100000;
				7'b0011101 : out = 8'b0011000;
				7'b0011110 : out = 8'b0010000;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0111001;
				7'b0100001 : out = 8'b0110001;
				7'b0100010 : out = 8'b0101001;
				7'b0100011 : out = 8'b0100001;
				7'b0100100 : out = 8'b0011001;
				7'b0100101 : out = 8'b0010001;
				7'b0100110 : out = 8'b0001001;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0111011;
				7'b0101001 : out = 8'b0110011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0100011;
				7'b0101100 : out = 8'b0011011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000011;
				7'b0110000 : out = 8'b0111101;
				7'b0110001 : out = 8'b0110101;
				7'b0110010 : out = 8'b0101101;
				7'b0110011 : out = 8'b0100101;
				7'b0110100 : out = 8'b0011101;
				7'b0110101 : out = 8'b0010101;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0000101;
				7'b0111000 : out = 8'b0111111;
				7'b0111001 : out = 8'b0110111;
				7'b0111010 : out = 8'b0101111;
				7'b0111011 : out = 8'b0100111;
				7'b0111100 : out = 8'b0011111;
				7'b0111101 : out = 8'b0010111;
				7'b0111110 : out = 8'b0001111;
				7'b0111111 : out = 8'b0000111;
			endcase
		  end

endmodule

module per(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b010000;
				6'b000001 : out = 8'b000111;
				6'b000010 : out = 8'b010100;
				6'b000011 : out = 8'b010101;
				6'b000100 : out = 8'b011101;
				6'b000101 : out = 8'b001100;
				6'b000110 : out = 8'b011100;
				6'b000111 : out = 8'b010001;
				6'b001000 : out = 8'b000001;
				6'b001001 : out = 8'b001111;
				6'b001010 : out = 8'b010111;
				6'b001011 : out = 8'b011010;
				6'b001100 : out = 8'b000101;
				6'b001101 : out = 8'b010010;
				6'b001110 : out = 8'b011111;
				6'b001111 : out = 8'b001010;
				6'b010000 : out = 8'b000010;
				6'b010001 : out = 8'b001000;
				6'b010010 : out = 8'b011000;
				6'b010011 : out = 8'b001110;
				6'b010100 : out = 8'b100000;
				6'b010101 : out = 8'b011011;
				6'b010110 : out = 8'b000011;
				6'b010111 : out = 8'b001001;
				6'b011000 : out = 8'b010011;
				6'b011001 : out = 8'b001101;
				6'b011010 : out = 8'b011110;
				6'b011011 : out = 8'b000110;
				6'b011100 : out = 8'b010110;
				6'b011101 : out = 8'b001011;
				6'b011110 : out = 8'b000100;
				6'b011111 : out = 8'b011001;
			endcase
		  end

endmodule

module sbox_0(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001110;
				7'b0000001 : out = 8'b0000100;
				7'b0000010 : out = 8'b0001101;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000010;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001010;
				7'b0001010 : out = 8'b0000110;
				7'b0001011 : out = 8'b0001100;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001001;
				7'b0001110 : out = 8'b0000000;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000000;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000111;
				7'b0010011 : out = 8'b0000100;
				7'b0010100 : out = 8'b0001110;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0001010;
				7'b0011001 : out = 8'b0000110;
				7'b0011010 : out = 8'b0001100;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0001001;
				7'b0011101 : out = 8'b0000101;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000001;
				7'b0100010 : out = 8'b0001110;
				7'b0100011 : out = 8'b0001000;
				7'b0100100 : out = 8'b0001101;
				7'b0100101 : out = 8'b0000110;
				7'b0100110 : out = 8'b0000010;
				7'b0100111 : out = 8'b0001011;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001100;
				7'b0101010 : out = 8'b0001001;
				7'b0101011 : out = 8'b0000111;
				7'b0101100 : out = 8'b0000011;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0000000;
				7'b0110000 : out = 8'b0001111;
				7'b0110001 : out = 8'b0001100;
				7'b0110010 : out = 8'b0001000;
				7'b0110011 : out = 8'b0000010;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0000001;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000101;
				7'b0111001 : out = 8'b0001011;
				7'b0111010 : out = 8'b0000011;
				7'b0111011 : out = 8'b0001110;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule

module sbox_1(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001111;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001011;
				7'b0000110 : out = 8'b0000011;
				7'b0000111 : out = 8'b0000100;
				7'b0001000 : out = 8'b0001001;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0000010;
				7'b0001011 : out = 8'b0001101;
				7'b0001100 : out = 8'b0001100;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001010;
				7'b0010000 : out = 8'b0000011;
				7'b0010001 : out = 8'b0001101;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0001111;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001000;
				7'b0010111 : out = 8'b0001110;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0000001;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000110;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001011;
				7'b0011111 : out = 8'b0000101;
				7'b0100000 : out = 8'b0000000;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0000111;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0000100;
				7'b0100110 : out = 8'b0001101;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0000101;
				7'b0101001 : out = 8'b0001000;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000110;
				7'b0101100 : out = 8'b0001001;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000010;
				7'b0101111 : out = 8'b0001111;
				7'b0110000 : out = 8'b0001101;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001010;
				7'b0110011 : out = 8'b0000001;
				7'b0110100 : out = 8'b0000011;
				7'b0110101 : out = 8'b0001111;
				7'b0110110 : out = 8'b0000100;
				7'b0110111 : out = 8'b0000010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0000110;
				7'b0111010 : out = 8'b0000111;
				7'b0111011 : out = 8'b0001100;
				7'b0111100 : out = 8'b0000000;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0001110;
				7'b0111111 : out = 8'b0001001;
			endcase
		  end

endmodule

module sbox_2(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001010;
				7'b0000001 : out = 8'b0000000;
				7'b0000010 : out = 8'b0001001;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0000011;
				7'b0000110 : out = 8'b0001111;
				7'b0000111 : out = 8'b0000101;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0001100;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0000100;
				7'b0001110 : out = 8'b0000010;
				7'b0001111 : out = 8'b0001000;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000111;
				7'b0010010 : out = 8'b0000000;
				7'b0010011 : out = 8'b0001001;
				7'b0010100 : out = 8'b0000011;
				7'b0010101 : out = 8'b0000100;
				7'b0010110 : out = 8'b0000110;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0000010;
				7'b0011001 : out = 8'b0001000;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0001100;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0001111;
				7'b0011111 : out = 8'b0000001;
				7'b0100000 : out = 8'b0001101;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0001001;
				7'b0100100 : out = 8'b0001000;
				7'b0100101 : out = 8'b0001111;
				7'b0100110 : out = 8'b0000011;
				7'b0100111 : out = 8'b0000000;
				7'b0101000 : out = 8'b0001011;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000010;
				7'b0101011 : out = 8'b0001100;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0001110;
				7'b0101111 : out = 8'b0000111;
				7'b0110000 : out = 8'b0000001;
				7'b0110001 : out = 8'b0001010;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0000000;
				7'b0110100 : out = 8'b0000110;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000100;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0001110;
				7'b0111011 : out = 8'b0000011;
				7'b0111100 : out = 8'b0001011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule

module sbox_3(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000111;
				7'b0000001 : out = 8'b0001101;
				7'b0000010 : out = 8'b0001110;
				7'b0000011 : out = 8'b0000011;
				7'b0000100 : out = 8'b0000000;
				7'b0000101 : out = 8'b0000110;
				7'b0000110 : out = 8'b0001001;
				7'b0000111 : out = 8'b0001010;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0000010;
				7'b0001010 : out = 8'b0001000;
				7'b0001011 : out = 8'b0000101;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0001100;
				7'b0001110 : out = 8'b0000100;
				7'b0001111 : out = 8'b0001111;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0001000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000101;
				7'b0010100 : out = 8'b0000110;
				7'b0010101 : out = 8'b0001111;
				7'b0010110 : out = 8'b0000000;
				7'b0010111 : out = 8'b0000011;
				7'b0011000 : out = 8'b0000100;
				7'b0011001 : out = 8'b0000111;
				7'b0011010 : out = 8'b0000010;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000001;
				7'b0011101 : out = 8'b0001010;
				7'b0011110 : out = 8'b0001110;
				7'b0011111 : out = 8'b0001001;
				7'b0100000 : out = 8'b0001010;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0001001;
				7'b0100011 : out = 8'b0000000;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0001011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001101;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000011;
				7'b0101011 : out = 8'b0001110;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0000010;
				7'b0101110 : out = 8'b0001000;
				7'b0101111 : out = 8'b0000100;
				7'b0110000 : out = 8'b0000011;
				7'b0110001 : out = 8'b0001111;
				7'b0110010 : out = 8'b0000000;
				7'b0110011 : out = 8'b0000110;
				7'b0110100 : out = 8'b0001010;
				7'b0110101 : out = 8'b0000001;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0001000;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000100;
				7'b0111010 : out = 8'b0000101;
				7'b0111011 : out = 8'b0001011;
				7'b0111100 : out = 8'b0001100;
				7'b0111101 : out = 8'b0000111;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001110;
			endcase
		  end

endmodule

module sbox_4(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000010;
				7'b0000001 : out = 8'b0001100;
				7'b0000010 : out = 8'b0000100;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000111;
				7'b0000101 : out = 8'b0001010;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000110;
				7'b0001000 : out = 8'b0001000;
				7'b0001001 : out = 8'b0000101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0001101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001110;
				7'b0001111 : out = 8'b0001001;
				7'b0010000 : out = 8'b0001110;
				7'b0010001 : out = 8'b0001011;
				7'b0010010 : out = 8'b0000010;
				7'b0010011 : out = 8'b0001100;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0000111;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0000101;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0001111;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000011;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000010;
				7'b0100010 : out = 8'b0000001;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0001101;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001000;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001001;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000101;
				7'b0101100 : out = 8'b0000110;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000000;
				7'b0101111 : out = 8'b0001110;
				7'b0110000 : out = 8'b0001011;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001100;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0001110;
				7'b0110110 : out = 8'b0000010;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0000110;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000100;
				7'b0111110 : out = 8'b0000101;
				7'b0111111 : out = 8'b0000011;
			endcase
		  end

endmodule

module sbox_5(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001100;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001010;
				7'b0000011 : out = 8'b0001111;
				7'b0000100 : out = 8'b0001001;
				7'b0000101 : out = 8'b0000010;
				7'b0000110 : out = 8'b0000110;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000000;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0000100;
				7'b0001100 : out = 8'b0001110;
				7'b0001101 : out = 8'b0000111;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001011;
				7'b0010000 : out = 8'b0001010;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000010;
				7'b0010100 : out = 8'b0000111;
				7'b0010101 : out = 8'b0001100;
				7'b0010110 : out = 8'b0001001;
				7'b0010111 : out = 8'b0000101;
				7'b0011000 : out = 8'b0000110;
				7'b0011001 : out = 8'b0000001;
				7'b0011010 : out = 8'b0001101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0001001;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0001111;
				7'b0100011 : out = 8'b0000101;
				7'b0100100 : out = 8'b0000010;
				7'b0100101 : out = 8'b0001000;
				7'b0100110 : out = 8'b0001100;
				7'b0100111 : out = 8'b0000011;
				7'b0101000 : out = 8'b0000111;
				7'b0101001 : out = 8'b0000000;
				7'b0101010 : out = 8'b0000100;
				7'b0101011 : out = 8'b0001010;
				7'b0101100 : out = 8'b0000001;
				7'b0101101 : out = 8'b0001101;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000110;
				7'b0110000 : out = 8'b0000100;
				7'b0110001 : out = 8'b0000011;
				7'b0110010 : out = 8'b0000010;
				7'b0110011 : out = 8'b0001100;
				7'b0110100 : out = 8'b0001001;
				7'b0110101 : out = 8'b0000101;
				7'b0110110 : out = 8'b0001111;
				7'b0110111 : out = 8'b0001010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0001110;
				7'b0111010 : out = 8'b0000001;
				7'b0111011 : out = 8'b0000111;
				7'b0111100 : out = 8'b0000110;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0001000;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule

module sbox_6(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000100;
				7'b0000001 : out = 8'b0001011;
				7'b0000010 : out = 8'b0000010;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0001111;
				7'b0000101 : out = 8'b0000000;
				7'b0000110 : out = 8'b0001000;
				7'b0000111 : out = 8'b0001101;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001100;
				7'b0001010 : out = 8'b0001001;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001010;
				7'b0001110 : out = 8'b0000110;
				7'b0001111 : out = 8'b0000001;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0001001;
				7'b0010110 : out = 8'b0000001;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0001110;
				7'b0011001 : out = 8'b0000011;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000010;
				7'b0011101 : out = 8'b0001111;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000001;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0001011;
				7'b0100011 : out = 8'b0001101;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0000011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001110;
				7'b0101000 : out = 8'b0001010;
				7'b0101001 : out = 8'b0001111;
				7'b0101010 : out = 8'b0000110;
				7'b0101011 : out = 8'b0001000;
				7'b0101100 : out = 8'b0000000;
				7'b0101101 : out = 8'b0000101;
				7'b0101110 : out = 8'b0001001;
				7'b0101111 : out = 8'b0000010;
				7'b0110000 : out = 8'b0000110;
				7'b0110001 : out = 8'b0001011;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0001000;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0000100;
				7'b0110110 : out = 8'b0001010;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000101;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001111;
				7'b0111100 : out = 8'b0001110;
				7'b0111101 : out = 8'b0000010;
				7'b0111110 : out = 8'b0000011;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule

module sbox_7(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001101;
				7'b0000001 : out = 8'b0000010;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0000100;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000001;
				7'b0001000 : out = 8'b0001010;
				7'b0001001 : out = 8'b0001001;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001110;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000001;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0001101;
				7'b0010011 : out = 8'b0001000;
				7'b0010100 : out = 8'b0001010;
				7'b0010101 : out = 8'b0000011;
				7'b0010110 : out = 8'b0000111;
				7'b0010111 : out = 8'b0000100;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0000110;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001110;
				7'b0011110 : out = 8'b0001001;
				7'b0011111 : out = 8'b0000010;
				7'b0100000 : out = 8'b0000111;
				7'b0100001 : out = 8'b0001011;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0000001;
				7'b0100100 : out = 8'b0001001;
				7'b0100101 : out = 8'b0001100;
				7'b0100110 : out = 8'b0001110;
				7'b0100111 : out = 8'b0000010;
				7'b0101000 : out = 8'b0000000;
				7'b0101001 : out = 8'b0000110;
				7'b0101010 : out = 8'b0001010;
				7'b0101011 : out = 8'b0001101;
				7'b0101100 : out = 8'b0001111;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0001000;
				7'b0110000 : out = 8'b0000010;
				7'b0110001 : out = 8'b0000001;
				7'b0110010 : out = 8'b0001110;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001010;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0001111;
				7'b0111001 : out = 8'b0001100;
				7'b0111010 : out = 8'b0001001;
				7'b0111011 : out = 8'b0000000;
				7'b0111100 : out = 8'b0000011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001011;
			endcase
		  end

endmodule

module exp_d(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b100000;
				6'b000001 : out = 8'b000001;
				6'b000010 : out = 8'b000010;
				6'b000011 : out = 8'b000011;
				6'b000100 : out = 8'b000100;
				6'b000101 : out = 8'b000101;
				6'b000110 : out = 8'b000100;
				6'b000111 : out = 8'b000101;
				6'b001000 : out = 8'b000110;
				6'b001001 : out = 8'b000111;
				6'b001010 : out = 8'b001000;
				6'b001011 : out = 8'b001001;
				6'b001100 : out = 8'b001000;
				6'b001101 : out = 8'b001001;
				6'b001110 : out = 8'b001010;
				6'b001111 : out = 8'b001011;
				6'b010000 : out = 8'b001100;
				6'b010001 : out = 8'b001101;
				6'b010010 : out = 8'b001100;
				6'b010011 : out = 8'b001101;
				6'b010100 : out = 8'b001110;
				6'b010101 : out = 8'b001111;
				6'b010110 : out = 8'b010000;
				6'b010111 : out = 8'b010001;
				6'b011000 : out = 8'b010000;
				6'b011001 : out = 8'b010001;
				6'b011010 : out = 8'b010010;
				6'b011011 : out = 8'b010011;
				6'b011100 : out = 8'b010100;
				6'b011101 : out = 8'b010101;
				6'b011110 : out = 8'b010100;
				6'b011111 : out = 8'b010101;
				6'b100000 : out = 8'b010110;
				6'b100001 : out = 8'b010111;
				6'b100010 : out = 8'b011000;
				6'b100011 : out = 8'b011001;
				6'b100100 : out = 8'b011000;
				6'b100101 : out = 8'b011001;
				6'b100110 : out = 8'b011010;
				6'b100111 : out = 8'b011011;
				6'b101000 : out = 8'b011100;
				6'b101001 : out = 8'b011101;
				6'b101010 : out = 8'b011100;
				6'b101011 : out = 8'b011101;
				6'b101100 : out = 8'b011110;
				6'b101101 : out = 8'b011111;
				6'b101110 : out = 8'b100000;
				6'b101111 : out = 8'b000001;
			endcase
		  end

endmodule


module final_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0101000;
				7'b0000001 : out = 8'b0001000;
				7'b0000010 : out = 8'b0110000;
				7'b0000011 : out = 8'b0010000;
				7'b0000100 : out = 8'b0111000;
				7'b0000101 : out = 8'b0011000;
				7'b0000110 : out = 8'b1000000;
				7'b0000111 : out = 8'b0100000;
				7'b0001000 : out = 8'b0100111;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0101111;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0110111;
				7'b0001101 : out = 8'b0010111;
				7'b0001110 : out = 8'b0111111;
				7'b0001111 : out = 8'b0011111;
				7'b0010000 : out = 8'b0100110;
				7'b0010001 : out = 8'b0000110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0001110;
				7'b0010100 : out = 8'b0110110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0111110;
				7'b0010111 : out = 8'b0011110;
				7'b0011000 : out = 8'b0100101;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0101101;
				7'b0011011 : out = 8'b0001101;
				7'b0011100 : out = 8'b0110101;
				7'b0011101 : out = 8'b0010101;
				7'b0011110 : out = 8'b0111101;
				7'b0011111 : out = 8'b0011101;
				7'b0100000 : out = 8'b0100100;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0101100;
				7'b0100011 : out = 8'b0001100;
				7'b0100100 : out = 8'b0110100;
				7'b0100101 : out = 8'b0010100;
				7'b0100110 : out = 8'b0111100;
				7'b0100111 : out = 8'b0011100;
				7'b0101000 : out = 8'b0100011;
				7'b0101001 : out = 8'b0000011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0001011;
				7'b0101100 : out = 8'b0110011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0111011;
				7'b0101111 : out = 8'b0011011;
				7'b0110000 : out = 8'b0100010;
				7'b0110001 : out = 8'b0000010;
				7'b0110010 : out = 8'b0101010;
				7'b0110011 : out = 8'b0001010;
				7'b0110100 : out = 8'b0110010;
				7'b0110101 : out = 8'b0010010;
				7'b0110110 : out = 8'b0111010;
				7'b0110111 : out = 8'b0011010;
				7'b0111000 : out = 8'b0100001;
				7'b0111001 : out = 8'b0000001;
				7'b0111010 : out = 8'b0101001;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0110001;
				7'b0111101 : out = 8'b0010001;
				7'b0111110 : out = 8'b0111001;
				7'b0111111 : out = 8'b0011001;
			endcase
		  end

endmodule


module initial_perm(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0111010;
				7'b0000001 : out = 8'b0110010;
				7'b0000010 : out = 8'b0101010;
				7'b0000011 : out = 8'b0100010;
				7'b0000100 : out = 8'b0011010;
				7'b0000101 : out = 8'b0010010;
				7'b0000110 : out = 8'b0001010;
				7'b0000111 : out = 8'b0000010;
				7'b0001000 : out = 8'b0111100;
				7'b0001001 : out = 8'b0110100;
				7'b0001010 : out = 8'b0101100;
				7'b0001011 : out = 8'b0100100;
				7'b0001100 : out = 8'b0011100;
				7'b0001101 : out = 8'b0010100;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000100;
				7'b0010000 : out = 8'b0111110;
				7'b0010001 : out = 8'b0110110;
				7'b0010010 : out = 8'b0101110;
				7'b0010011 : out = 8'b0100110;
				7'b0010100 : out = 8'b0011110;
				7'b0010101 : out = 8'b0010110;
				7'b0010110 : out = 8'b0001110;
				7'b0010111 : out = 8'b0000110;
				7'b0011000 : out = 8'b1000000;
				7'b0011001 : out = 8'b0111000;
				7'b0011010 : out = 8'b0110000;
				7'b0011011 : out = 8'b0101000;
				7'b0011100 : out = 8'b0100000;
				7'b0011101 : out = 8'b0011000;
				7'b0011110 : out = 8'b0010000;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0111001;
				7'b0100001 : out = 8'b0110001;
				7'b0100010 : out = 8'b0101001;
				7'b0100011 : out = 8'b0100001;
				7'b0100100 : out = 8'b0011001;
				7'b0100101 : out = 8'b0010001;
				7'b0100110 : out = 8'b0001001;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0111011;
				7'b0101001 : out = 8'b0110011;
				7'b0101010 : out = 8'b0101011;
				7'b0101011 : out = 8'b0100011;
				7'b0101100 : out = 8'b0011011;
				7'b0101101 : out = 8'b0010011;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000011;
				7'b0110000 : out = 8'b0111101;
				7'b0110001 : out = 8'b0110101;
				7'b0110010 : out = 8'b0101101;
				7'b0110011 : out = 8'b0100101;
				7'b0110100 : out = 8'b0011101;
				7'b0110101 : out = 8'b0010101;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0000101;
				7'b0111000 : out = 8'b0111111;
				7'b0111001 : out = 8'b0110111;
				7'b0111010 : out = 8'b0101111;
				7'b0111011 : out = 8'b0100111;
				7'b0111100 : out = 8'b0011111;
				7'b0111101 : out = 8'b0010111;
				7'b0111110 : out = 8'b0001111;
				7'b0111111 : out = 8'b0000111;
			endcase
		  end

endmodule


module per(input logic [5:0] in,
		output logic [5:0] out);

		always_comb
		  begin
			case(in)
				6'b000000 : out = 8'b010000;
				6'b000001 : out = 8'b000111;
				6'b000010 : out = 8'b010100;
				6'b000011 : out = 8'b010101;
				6'b000100 : out = 8'b011101;
				6'b000101 : out = 8'b001100;
				6'b000110 : out = 8'b011100;
				6'b000111 : out = 8'b010001;
				6'b001000 : out = 8'b000001;
				6'b001001 : out = 8'b001111;
				6'b001010 : out = 8'b010111;
				6'b001011 : out = 8'b011010;
				6'b001100 : out = 8'b000101;
				6'b001101 : out = 8'b010010;
				6'b001110 : out = 8'b011111;
				6'b001111 : out = 8'b001010;
				6'b010000 : out = 8'b000010;
				6'b010001 : out = 8'b001000;
				6'b010010 : out = 8'b011000;
				6'b010011 : out = 8'b001110;
				6'b010100 : out = 8'b100000;
				6'b010101 : out = 8'b011011;
				6'b010110 : out = 8'b000011;
				6'b010111 : out = 8'b001001;
				6'b011000 : out = 8'b010011;
				6'b011001 : out = 8'b001101;
				6'b011010 : out = 8'b011110;
				6'b011011 : out = 8'b000110;
				6'b011100 : out = 8'b010110;
				6'b011101 : out = 8'b001011;
				6'b011110 : out = 8'b000100;
				6'b011111 : out = 8'b011001;
			endcase
		  end

endmodule


module sbox_0(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001110;
				7'b0000001 : out = 8'b0000100;
				7'b0000010 : out = 8'b0001101;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000010;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001010;
				7'b0001010 : out = 8'b0000110;
				7'b0001011 : out = 8'b0001100;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001001;
				7'b0001110 : out = 8'b0000000;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000000;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000111;
				7'b0010011 : out = 8'b0000100;
				7'b0010100 : out = 8'b0001110;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0001010;
				7'b0011001 : out = 8'b0000110;
				7'b0011010 : out = 8'b0001100;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0001001;
				7'b0011101 : out = 8'b0000101;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000001;
				7'b0100010 : out = 8'b0001110;
				7'b0100011 : out = 8'b0001000;
				7'b0100100 : out = 8'b0001101;
				7'b0100101 : out = 8'b0000110;
				7'b0100110 : out = 8'b0000010;
				7'b0100111 : out = 8'b0001011;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001100;
				7'b0101010 : out = 8'b0001001;
				7'b0101011 : out = 8'b0000111;
				7'b0101100 : out = 8'b0000011;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0000000;
				7'b0110000 : out = 8'b0001111;
				7'b0110001 : out = 8'b0001100;
				7'b0110010 : out = 8'b0001000;
				7'b0110011 : out = 8'b0000010;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0000001;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000101;
				7'b0111001 : out = 8'b0001011;
				7'b0111010 : out = 8'b0000011;
				7'b0111011 : out = 8'b0001110;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule


module sbox_1(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001111;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001011;
				7'b0000110 : out = 8'b0000011;
				7'b0000111 : out = 8'b0000100;
				7'b0001000 : out = 8'b0001001;
				7'b0001001 : out = 8'b0000111;
				7'b0001010 : out = 8'b0000010;
				7'b0001011 : out = 8'b0001101;
				7'b0001100 : out = 8'b0001100;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001010;
				7'b0010000 : out = 8'b0000011;
				7'b0010001 : out = 8'b0001101;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0001111;
				7'b0010101 : out = 8'b0000010;
				7'b0010110 : out = 8'b0001000;
				7'b0010111 : out = 8'b0001110;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0000001;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000110;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001011;
				7'b0011111 : out = 8'b0000101;
				7'b0100000 : out = 8'b0000000;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0000111;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0000100;
				7'b0100110 : out = 8'b0001101;
				7'b0100111 : out = 8'b0000001;
				7'b0101000 : out = 8'b0000101;
				7'b0101001 : out = 8'b0001000;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000110;
				7'b0101100 : out = 8'b0001001;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000010;
				7'b0101111 : out = 8'b0001111;
				7'b0110000 : out = 8'b0001101;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001010;
				7'b0110011 : out = 8'b0000001;
				7'b0110100 : out = 8'b0000011;
				7'b0110101 : out = 8'b0001111;
				7'b0110110 : out = 8'b0000100;
				7'b0110111 : out = 8'b0000010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0000110;
				7'b0111010 : out = 8'b0000111;
				7'b0111011 : out = 8'b0001100;
				7'b0111100 : out = 8'b0000000;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0001110;
				7'b0111111 : out = 8'b0001001;
			endcase
		  end

endmodule


module sbox_2(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001010;
				7'b0000001 : out = 8'b0000000;
				7'b0000010 : out = 8'b0001001;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0000011;
				7'b0000110 : out = 8'b0001111;
				7'b0000111 : out = 8'b0000101;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0001100;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0000100;
				7'b0001110 : out = 8'b0000010;
				7'b0001111 : out = 8'b0001000;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000111;
				7'b0010010 : out = 8'b0000000;
				7'b0010011 : out = 8'b0001001;
				7'b0010100 : out = 8'b0000011;
				7'b0010101 : out = 8'b0000100;
				7'b0010110 : out = 8'b0000110;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0000010;
				7'b0011001 : out = 8'b0001000;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0001100;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0001111;
				7'b0011111 : out = 8'b0000001;
				7'b0100000 : out = 8'b0001101;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0001001;
				7'b0100100 : out = 8'b0001000;
				7'b0100101 : out = 8'b0001111;
				7'b0100110 : out = 8'b0000011;
				7'b0100111 : out = 8'b0000000;
				7'b0101000 : out = 8'b0001011;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000010;
				7'b0101011 : out = 8'b0001100;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0001010;
				7'b0101110 : out = 8'b0001110;
				7'b0101111 : out = 8'b0000111;
				7'b0110000 : out = 8'b0000001;
				7'b0110001 : out = 8'b0001010;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0000000;
				7'b0110100 : out = 8'b0000110;
				7'b0110101 : out = 8'b0001001;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0000100;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0001110;
				7'b0111011 : out = 8'b0000011;
				7'b0111100 : out = 8'b0001011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule


module sbox_3(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000111;
				7'b0000001 : out = 8'b0001101;
				7'b0000010 : out = 8'b0001110;
				7'b0000011 : out = 8'b0000011;
				7'b0000100 : out = 8'b0000000;
				7'b0000101 : out = 8'b0000110;
				7'b0000110 : out = 8'b0001001;
				7'b0000111 : out = 8'b0001010;
				7'b0001000 : out = 8'b0000001;
				7'b0001001 : out = 8'b0000010;
				7'b0001010 : out = 8'b0001000;
				7'b0001011 : out = 8'b0000101;
				7'b0001100 : out = 8'b0001011;
				7'b0001101 : out = 8'b0001100;
				7'b0001110 : out = 8'b0000100;
				7'b0001111 : out = 8'b0001111;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0001000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000101;
				7'b0010100 : out = 8'b0000110;
				7'b0010101 : out = 8'b0001111;
				7'b0010110 : out = 8'b0000000;
				7'b0010111 : out = 8'b0000011;
				7'b0011000 : out = 8'b0000100;
				7'b0011001 : out = 8'b0000111;
				7'b0011010 : out = 8'b0000010;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000001;
				7'b0011101 : out = 8'b0001010;
				7'b0011110 : out = 8'b0001110;
				7'b0011111 : out = 8'b0001001;
				7'b0100000 : out = 8'b0001010;
				7'b0100001 : out = 8'b0000110;
				7'b0100010 : out = 8'b0001001;
				7'b0100011 : out = 8'b0000000;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0001011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001101;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0000001;
				7'b0101010 : out = 8'b0000011;
				7'b0101011 : out = 8'b0001110;
				7'b0101100 : out = 8'b0000101;
				7'b0101101 : out = 8'b0000010;
				7'b0101110 : out = 8'b0001000;
				7'b0101111 : out = 8'b0000100;
				7'b0110000 : out = 8'b0000011;
				7'b0110001 : out = 8'b0001111;
				7'b0110010 : out = 8'b0000000;
				7'b0110011 : out = 8'b0000110;
				7'b0110100 : out = 8'b0001010;
				7'b0110101 : out = 8'b0000001;
				7'b0110110 : out = 8'b0001101;
				7'b0110111 : out = 8'b0001000;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000100;
				7'b0111010 : out = 8'b0000101;
				7'b0111011 : out = 8'b0001011;
				7'b0111100 : out = 8'b0001100;
				7'b0111101 : out = 8'b0000111;
				7'b0111110 : out = 8'b0000010;
				7'b0111111 : out = 8'b0001110;
			endcase
		  end

endmodule


module sbox_4(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000010;
				7'b0000001 : out = 8'b0001100;
				7'b0000010 : out = 8'b0000100;
				7'b0000011 : out = 8'b0000001;
				7'b0000100 : out = 8'b0000111;
				7'b0000101 : out = 8'b0001010;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000110;
				7'b0001000 : out = 8'b0001000;
				7'b0001001 : out = 8'b0000101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001111;
				7'b0001100 : out = 8'b0001101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001110;
				7'b0001111 : out = 8'b0001001;
				7'b0010000 : out = 8'b0001110;
				7'b0010001 : out = 8'b0001011;
				7'b0010010 : out = 8'b0000010;
				7'b0010011 : out = 8'b0001100;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0000111;
				7'b0010110 : out = 8'b0001101;
				7'b0010111 : out = 8'b0000001;
				7'b0011000 : out = 8'b0000101;
				7'b0011001 : out = 8'b0000000;
				7'b0011010 : out = 8'b0001111;
				7'b0011011 : out = 8'b0001010;
				7'b0011100 : out = 8'b0000011;
				7'b0011101 : out = 8'b0001001;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000100;
				7'b0100001 : out = 8'b0000010;
				7'b0100010 : out = 8'b0000001;
				7'b0100011 : out = 8'b0001011;
				7'b0100100 : out = 8'b0001010;
				7'b0100101 : out = 8'b0001101;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001000;
				7'b0101000 : out = 8'b0001111;
				7'b0101001 : out = 8'b0001001;
				7'b0101010 : out = 8'b0001100;
				7'b0101011 : out = 8'b0000101;
				7'b0101100 : out = 8'b0000110;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000000;
				7'b0101111 : out = 8'b0001110;
				7'b0110000 : out = 8'b0001011;
				7'b0110001 : out = 8'b0001000;
				7'b0110010 : out = 8'b0001100;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0001110;
				7'b0110110 : out = 8'b0000010;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0000110;
				7'b0111001 : out = 8'b0001111;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001001;
				7'b0111100 : out = 8'b0001010;
				7'b0111101 : out = 8'b0000100;
				7'b0111110 : out = 8'b0000101;
				7'b0111111 : out = 8'b0000011;
			endcase
		  end

endmodule


module sbox_5(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001100;
				7'b0000001 : out = 8'b0000001;
				7'b0000010 : out = 8'b0001010;
				7'b0000011 : out = 8'b0001111;
				7'b0000100 : out = 8'b0001001;
				7'b0000101 : out = 8'b0000010;
				7'b0000110 : out = 8'b0000110;
				7'b0000111 : out = 8'b0001000;
				7'b0001000 : out = 8'b0000000;
				7'b0001001 : out = 8'b0001101;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0000100;
				7'b0001100 : out = 8'b0001110;
				7'b0001101 : out = 8'b0000111;
				7'b0001110 : out = 8'b0000101;
				7'b0001111 : out = 8'b0001011;
				7'b0010000 : out = 8'b0001010;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0000100;
				7'b0010011 : out = 8'b0000010;
				7'b0010100 : out = 8'b0000111;
				7'b0010101 : out = 8'b0001100;
				7'b0010110 : out = 8'b0001001;
				7'b0010111 : out = 8'b0000101;
				7'b0011000 : out = 8'b0000110;
				7'b0011001 : out = 8'b0000001;
				7'b0011010 : out = 8'b0001101;
				7'b0011011 : out = 8'b0001110;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001011;
				7'b0011110 : out = 8'b0000011;
				7'b0011111 : out = 8'b0001000;
				7'b0100000 : out = 8'b0001001;
				7'b0100001 : out = 8'b0001110;
				7'b0100010 : out = 8'b0001111;
				7'b0100011 : out = 8'b0000101;
				7'b0100100 : out = 8'b0000010;
				7'b0100101 : out = 8'b0001000;
				7'b0100110 : out = 8'b0001100;
				7'b0100111 : out = 8'b0000011;
				7'b0101000 : out = 8'b0000111;
				7'b0101001 : out = 8'b0000000;
				7'b0101010 : out = 8'b0000100;
				7'b0101011 : out = 8'b0001010;
				7'b0101100 : out = 8'b0000001;
				7'b0101101 : out = 8'b0001101;
				7'b0101110 : out = 8'b0001011;
				7'b0101111 : out = 8'b0000110;
				7'b0110000 : out = 8'b0000100;
				7'b0110001 : out = 8'b0000011;
				7'b0110010 : out = 8'b0000010;
				7'b0110011 : out = 8'b0001100;
				7'b0110100 : out = 8'b0001001;
				7'b0110101 : out = 8'b0000101;
				7'b0110110 : out = 8'b0001111;
				7'b0110111 : out = 8'b0001010;
				7'b0111000 : out = 8'b0001011;
				7'b0111001 : out = 8'b0001110;
				7'b0111010 : out = 8'b0000001;
				7'b0111011 : out = 8'b0000111;
				7'b0111100 : out = 8'b0000110;
				7'b0111101 : out = 8'b0000000;
				7'b0111110 : out = 8'b0001000;
				7'b0111111 : out = 8'b0001101;
			endcase
		  end

endmodule


module sbox_6(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0000100;
				7'b0000001 : out = 8'b0001011;
				7'b0000010 : out = 8'b0000010;
				7'b0000011 : out = 8'b0001110;
				7'b0000100 : out = 8'b0001111;
				7'b0000101 : out = 8'b0000000;
				7'b0000110 : out = 8'b0001000;
				7'b0000111 : out = 8'b0001101;
				7'b0001000 : out = 8'b0000011;
				7'b0001001 : out = 8'b0001100;
				7'b0001010 : out = 8'b0001001;
				7'b0001011 : out = 8'b0000111;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0001010;
				7'b0001110 : out = 8'b0000110;
				7'b0001111 : out = 8'b0000001;
				7'b0010000 : out = 8'b0001101;
				7'b0010001 : out = 8'b0000000;
				7'b0010010 : out = 8'b0001011;
				7'b0010011 : out = 8'b0000111;
				7'b0010100 : out = 8'b0000100;
				7'b0010101 : out = 8'b0001001;
				7'b0010110 : out = 8'b0000001;
				7'b0010111 : out = 8'b0001010;
				7'b0011000 : out = 8'b0001110;
				7'b0011001 : out = 8'b0000011;
				7'b0011010 : out = 8'b0000101;
				7'b0011011 : out = 8'b0001100;
				7'b0011100 : out = 8'b0000010;
				7'b0011101 : out = 8'b0001111;
				7'b0011110 : out = 8'b0001000;
				7'b0011111 : out = 8'b0000110;
				7'b0100000 : out = 8'b0000001;
				7'b0100001 : out = 8'b0000100;
				7'b0100010 : out = 8'b0001011;
				7'b0100011 : out = 8'b0001101;
				7'b0100100 : out = 8'b0001100;
				7'b0100101 : out = 8'b0000011;
				7'b0100110 : out = 8'b0000111;
				7'b0100111 : out = 8'b0001110;
				7'b0101000 : out = 8'b0001010;
				7'b0101001 : out = 8'b0001111;
				7'b0101010 : out = 8'b0000110;
				7'b0101011 : out = 8'b0001000;
				7'b0101100 : out = 8'b0000000;
				7'b0101101 : out = 8'b0000101;
				7'b0101110 : out = 8'b0001001;
				7'b0101111 : out = 8'b0000010;
				7'b0110000 : out = 8'b0000110;
				7'b0110001 : out = 8'b0001011;
				7'b0110010 : out = 8'b0001101;
				7'b0110011 : out = 8'b0001000;
				7'b0110100 : out = 8'b0000001;
				7'b0110101 : out = 8'b0000100;
				7'b0110110 : out = 8'b0001010;
				7'b0110111 : out = 8'b0000111;
				7'b0111000 : out = 8'b0001001;
				7'b0111001 : out = 8'b0000101;
				7'b0111010 : out = 8'b0000000;
				7'b0111011 : out = 8'b0001111;
				7'b0111100 : out = 8'b0001110;
				7'b0111101 : out = 8'b0000010;
				7'b0111110 : out = 8'b0000011;
				7'b0111111 : out = 8'b0001100;
			endcase
		  end

endmodule


module sbox_7(input logic [6:0] in,
		output logic [6:0] out);

		always_comb
		  begin
			case(in)
				7'b0000000 : out = 8'b0001101;
				7'b0000001 : out = 8'b0000010;
				7'b0000010 : out = 8'b0001000;
				7'b0000011 : out = 8'b0000100;
				7'b0000100 : out = 8'b0000110;
				7'b0000101 : out = 8'b0001111;
				7'b0000110 : out = 8'b0001011;
				7'b0000111 : out = 8'b0000001;
				7'b0001000 : out = 8'b0001010;
				7'b0001001 : out = 8'b0001001;
				7'b0001010 : out = 8'b0000011;
				7'b0001011 : out = 8'b0001110;
				7'b0001100 : out = 8'b0000101;
				7'b0001101 : out = 8'b0000000;
				7'b0001110 : out = 8'b0001100;
				7'b0001111 : out = 8'b0000111;
				7'b0010000 : out = 8'b0000001;
				7'b0010001 : out = 8'b0001111;
				7'b0010010 : out = 8'b0001101;
				7'b0010011 : out = 8'b0001000;
				7'b0010100 : out = 8'b0001010;
				7'b0010101 : out = 8'b0000011;
				7'b0010110 : out = 8'b0000111;
				7'b0010111 : out = 8'b0000100;
				7'b0011000 : out = 8'b0001100;
				7'b0011001 : out = 8'b0000101;
				7'b0011010 : out = 8'b0000110;
				7'b0011011 : out = 8'b0001011;
				7'b0011100 : out = 8'b0000000;
				7'b0011101 : out = 8'b0001110;
				7'b0011110 : out = 8'b0001001;
				7'b0011111 : out = 8'b0000010;
				7'b0100000 : out = 8'b0000111;
				7'b0100001 : out = 8'b0001011;
				7'b0100010 : out = 8'b0000100;
				7'b0100011 : out = 8'b0000001;
				7'b0100100 : out = 8'b0001001;
				7'b0100101 : out = 8'b0001100;
				7'b0100110 : out = 8'b0001110;
				7'b0100111 : out = 8'b0000010;
				7'b0101000 : out = 8'b0000000;
				7'b0101001 : out = 8'b0000110;
				7'b0101010 : out = 8'b0001010;
				7'b0101011 : out = 8'b0001101;
				7'b0101100 : out = 8'b0001111;
				7'b0101101 : out = 8'b0000011;
				7'b0101110 : out = 8'b0000101;
				7'b0101111 : out = 8'b0001000;
				7'b0110000 : out = 8'b0000010;
				7'b0110001 : out = 8'b0000001;
				7'b0110010 : out = 8'b0001110;
				7'b0110011 : out = 8'b0000111;
				7'b0110100 : out = 8'b0000100;
				7'b0110101 : out = 8'b0001010;
				7'b0110110 : out = 8'b0001000;
				7'b0110111 : out = 8'b0001101;
				7'b0111000 : out = 8'b0001111;
				7'b0111001 : out = 8'b0001100;
				7'b0111010 : out = 8'b0001001;
				7'b0111011 : out = 8'b0000000;
				7'b0111100 : out = 8'b0000011;
				7'b0111101 : out = 8'b0000101;
				7'b0111110 : out = 8'b0000110;
				7'b0111111 : out = 8'b0001011;
			endcase
		  end

endmodule



/*
 Data Encryption Standard (S-DES)
 64-bit 16-round block cipher encryption and decryption algorithm 
 using 56-bit key (64-bit key with Parity).
 */

module GenerateKeys (Key, SubKey1, SubKey2, SubKey3, SubKey4,
		     SubKey5, SubKey6, SubKey7, SubKey8,
		     SubKey9, SubKey10, SubKey11, SubKey12,
		     SubKey13, SubKey14, SubKey15, SubKey16);
   
   // Generate SubKeys
   input logic [63:0]  Key;
   output logic [47:0] SubKey1;
   output logic [47:0] SubKey2;
   output logic [47:0] SubKey3;
   output logic [47:0] SubKey4;
   output logic [47:0] SubKey5;
   output logic [47:0] SubKey6;
   output logic [47:0] SubKey7;
   output logic [47:0] SubKey8;
   output logic [47:0] SubKey9;
   output logic [47:0] SubKey10;
   output logic [47:0] SubKey11;
   output logic [47:0] SubKey12;
   output logic [47:0] SubKey13;
   output logic [47:0] SubKey14;
   output logic [47:0] SubKey15;
   output logic [47:0] SubKey16;

   logic [27:0]        left_block0, left_block1, left_block2, left_block3;
   logic [27:0]        left_block4, left_block5, left_block6, left_block7;
   logic [27:0]        left_block8, left_block9, left_block10, left_block11;
   logic [27:0]        left_block12, left_block13, left_block14, left_block15;
   logic [27:0]        left_block16;
   logic [27:0]        right_block0, right_block1, right_block2, right_block3;
   logic [27:0]        right_block4, right_block5, right_block6, right_block7;
   logic [27:0]        right_block8, right_block9, right_block10, right_block11;
   logic [27:0]        right_block12, right_block13, right_block14, right_block15;
   logic [27:0]        right_block16;

   // Permutation Choice
   PC1 b1 (Key, left_block0, right_block0);

   // Perform each subkey using Rotate/Permutation Choice 2 (PC-2)
   // subkey 1      
   assign left_block1 = {left_block0[26:0], left_block0[27]};
   assign right_block1 = {right_block0[26:0], right_block0[27]};
   PC2 b2 (left_block1, right_block1, SubKey1);
   // subkey 2      
   assign left_block2 = {left_block1[26:0], left_block1[27]};
   assign right_block2 = {right_block1[26:0], right_block1[27]};
   PC2 b3 (left_block2, right_block2, SubKey2);
   // subkey 3
   assign left_block3 = {left_block2[25:0], left_block2[27:26]};
   assign right_block3 = {right_block2[25:0], right_block2[27:26]};
   PC2 b4 (left_block3, right_block3, SubKey3);
   // subkey 4
   assign left_block4 = {left_block3[25:0], left_block3[27:26]};
   assign right_block4 = {right_block3[25:0], right_block3[27:26]};
   PC2 b5 (left_block4, right_block4, SubKey4);
   // subkey 5
   assign left_block5 = {left_block4[25:0], left_block4[27:26]};
   assign right_block5 = {right_block4[25:0], right_block4[27:26]};
   PC2 b6 (left_block5, right_block5, SubKey5);
   // subkey 6
   assign left_block6 = {left_block5[25:0], left_block5[27:26]};
   assign right_block6 = {right_block5[25:0], right_block5[27:26]};
   PC2 b7 (left_block6, right_block6, SubKey6);
   // subkey 7
   assign left_block7 = {left_block6[25:0], left_block6[27:26]};
   assign right_block7 = {right_block6[25:0], right_block6[27:26]};
   PC2 b8 (left_block7, right_block7, SubKey7);
   // subkey 8
   assign left_block8 = {left_block7[25:0], left_block7[27:26]};
   assign right_block8 = {right_block7[25:0], right_block7[27:26]};
   PC2 b9 (left_block8, right_block8, SubKey8);                  
   // subkey 9      
   assign left_block9 = {left_block8[26:0], left_block8[27]};
   assign right_block9 = {right_block8[26:0], right_block8[27]};
   PC2 b10 (left_block9, right_block9, SubKey9);
   // subkey 10      
   assign left_block10 = {left_block9[25:0], left_block9[27:26]};
   assign right_block10 = {right_block9[25:0], right_block9[27:26]};
   PC2 b11 (left_block10, right_block10, SubKey10);
   // subkey 11     
   assign left_block11 = {left_block10[25:0], left_block10[27:26]};
   assign right_block11 = {right_block10[25:0], right_block10[27:26]};
   PC2 b12 (left_block11, right_block11, SubKey11);
   // subkey 12
   assign left_block12 = {left_block11[25:0], left_block11[27:26]};
   assign right_block12 = {right_block11[25:0], right_block11[27:26]};
   PC2 b13 (left_block12, right_block12, SubKey12);
   // subkey 13
   assign left_block13 = {left_block12[25:0], left_block12[27:26]};
   assign right_block13 = {right_block12[25:0], right_block12[27:26]};
   PC2 b14 (left_block13, right_block13, SubKey13);
   // subkey 14
   assign left_block14 = {left_block13[25:0], left_block13[27:26]};
   assign right_block14 = {right_block13[25:0], right_block13[27:26]};
   PC2 b15 (left_block14, right_block14, SubKey14);
   // subkey 15
   assign left_block15 = {left_block14[25:0], left_block14[27:26]};
   assign right_block15 = {right_block14[25:0], right_block14[27:26]};
   PC2 b16 (left_block15, right_block15, SubKey15);
   // subkey 16
   assign left_block16 = {left_block15[26:0], left_block15[27]};
   assign right_block16 = {right_block15[26:0], right_block15[27]};
   PC2 b17 (left_block16, right_block16, SubKey16);
   
endmodule // GenerateKeys

module PC1 (key, left_block, right_block);

   input logic [63:0]  key;
   output logic [27:0] left_block;
   output logic [27:0] right_block;

   logic [55:0]        out_block;

   assign {left_block, right_block} = out_block;
	
   assign out_block[55] = key[64-57];
   assign out_block[54] = key[64-49];
   assign out_block[53] = key[64-41];
   assign out_block[52] = key[64-33];
   assign out_block[51] = key[64-25];
   assign out_block[50] = key[64-17];
   assign out_block[49] = key[64-9];
   assign out_block[48] = key[64-1];
   assign out_block[47] = key[64-58];
   assign out_block[46] = key[64-50];
   assign out_block[45] = key[64-42];
   assign out_block[44] = key[64-34];
   assign out_block[43] = key[64-26];
   assign out_block[42] = key[64-18];
   assign out_block[41] = key[64-10];
   assign out_block[40] = key[64-2];
   assign out_block[39] = key[64-59];
   assign out_block[38] = key[64-51];
   assign out_block[37] = key[64-43];
   assign out_block[36] = key[64-35];
   assign out_block[35] = key[64-27];
   assign out_block[34] = key[64-19];
   assign out_block[33] = key[64-11];
   assign out_block[32] = key[64-3];
   assign out_block[31] = key[64-60];
   assign out_block[30] = key[64-52];
   assign out_block[29] = key[64-44];
   assign out_block[28] = key[64-36];
   assign out_block[27] = key[64-63];
   assign out_block[26] = key[64-55];
   assign out_block[25] = key[64-47];
   assign out_block[24] = key[64-39];
   assign out_block[23] = key[64-31];
   assign out_block[22] = key[64-23];
   assign out_block[21] = key[64-15];
   assign out_block[20] = key[64-7];
   assign out_block[19] = key[64-62];
   assign out_block[18] = key[64-54];
   assign out_block[17] = key[64-46];
   assign out_block[16] = key[64-38];
   assign out_block[15] = key[64-30];
   assign out_block[14] = key[64-22];
   assign out_block[13] = key[64-14];
   assign out_block[12] = key[64-6];
   assign out_block[11] = key[64-61];
   assign out_block[10] = key[64-53];
   assign out_block[9] = key[64-45];
   assign out_block[8] = key[64-37];
   assign out_block[7] = key[64-29];
   assign out_block[6] = key[64-21];
   assign out_block[5] = key[64-13];
   assign out_block[4] = key[64-5];
   assign out_block[3] = key[64-28];
   assign out_block[2] = key[64-20];
   assign out_block[1] = key[64-12];
   assign out_block[0] = key[64-4];

endmodule // PC1

module PC2 (left_block, right_block, subkey);

   input logic [27:0] left_block;
   input logic [27:0] right_block;
   output logic [47:0] subkey;

   logic [55:0]        combined;   

   assign combined = {left_block, right_block};
   
   assign subkey[47] = combined[56-14];
   assign subkey[46] = combined[56-17];
   assign subkey[45] = combined[56-11];
   assign subkey[44] = combined[56-24];
   assign subkey[43] = combined[56-1];
   assign subkey[42] = combined[56-5];
   assign subkey[41] = combined[56-3];
   assign subkey[40] = combined[56-28];
   assign subkey[39] = combined[56-15];
   assign subkey[38] = combined[56-6];   
   assign subkey[37] = combined[56-21];
   assign subkey[36] = combined[56-10];
   assign subkey[35] = combined[56-23];
   assign subkey[34] = combined[56-19];
   assign subkey[33] = combined[56-12];
   assign subkey[32] = combined[56-4];
   assign subkey[31] = combined[56-26];
   assign subkey[30] = combined[56-8];
   assign subkey[29] = combined[56-16];
   assign subkey[28] = combined[56-7];   
   assign subkey[27] = combined[56-27];
   assign subkey[26] = combined[56-20];
   assign subkey[25] = combined[56-13];
   assign subkey[24] = combined[56-2];
   assign subkey[23] = combined[56-41];
   assign subkey[22] = combined[56-52];
   assign subkey[21] = combined[56-31];
   assign subkey[20] = combined[56-37];
   assign subkey[19] = combined[56-47];
   assign subkey[18] = combined[56-55];   
   assign subkey[17] = combined[56-30];
   assign subkey[16] = combined[56-40];
   assign subkey[15] = combined[56-51];
   assign subkey[14] = combined[56-45];
   assign subkey[13] = combined[56-33];
   assign subkey[12] = combined[56-48];
   assign subkey[11] = combined[56-44];
   assign subkey[10] = combined[56-49];
   assign subkey[9] = combined[56-39];
   assign subkey[8] = combined[56-56];   
   assign subkey[7] = combined[56-34];
   assign subkey[6] = combined[56-53];
   assign subkey[5] = combined[56-46];
   assign subkey[4] = combined[56-42];
   assign subkey[3] = combined[56-50];
   assign subkey[2] = combined[56-36];
   assign subkey[1] = combined[56-29];
   assign subkey[0] = combined[56-32];
   
endmodule // PC2

// Straight Function
module SF (inp_block, out_block);

   input logic [31:0] inp_block;
   output logic [31:0] out_block;

   assign out_block[31] = inp_block[32-16];
   assign out_block[30] = inp_block[32-7];
   assign out_block[29] = inp_block[32-20];
   assign out_block[28] = inp_block[32-21];   
   assign out_block[27] = inp_block[32-29];
   assign out_block[26] = inp_block[32-12];
   assign out_block[25] = inp_block[32-28];
   assign out_block[24] = inp_block[32-17];
   assign out_block[23] = inp_block[32-1];
   assign out_block[22] = inp_block[32-15];
   assign out_block[21] = inp_block[32-23];
   assign out_block[20] = inp_block[32-26];
   assign out_block[19] = inp_block[32-5];
   assign out_block[18] = inp_block[32-18];   
   assign out_block[17] = inp_block[32-31];
   assign out_block[16] = inp_block[32-10];
   assign out_block[15] = inp_block[32-2];
   assign out_block[14] = inp_block[32-8];
   assign out_block[13] = inp_block[32-24];
   assign out_block[12] = inp_block[32-14];
   assign out_block[11] = inp_block[32-32];
   assign out_block[10] = inp_block[32-27];
   assign out_block[9] = inp_block[32-3];
   assign out_block[8] = inp_block[32-9];   
   assign out_block[7] = inp_block[32-19];
   assign out_block[6] = inp_block[32-13];
   assign out_block[5] = inp_block[32-30];
   assign out_block[4] = inp_block[32-6];
   assign out_block[3] = inp_block[32-22];
   assign out_block[2] = inp_block[32-11];
   assign out_block[1] = inp_block[32-4];
   assign out_block[0] = inp_block[32-25];

/* -----\/----- EXCLUDED -----\/-----
   assign out_block[ 0] = inp_block[16-1];
   assign out_block[ 1] = inp_block[7-1 ];
   assign out_block[ 2] = inp_block[20-1];
   assign out_block[ 3] = inp_block[21-1];   
   assign out_block[ 4] = inp_block[29-1];
   assign out_block[ 5] = inp_block[12-1];
   assign out_block[ 6] = inp_block[28-1];
   assign out_block[ 7] = inp_block[17-1];
   assign out_block[ 8] = inp_block[1-1 ];
   assign out_block[ 9] = inp_block[15-1];
   assign out_block[10] = inp_block[23-1];
   assign out_block[11] = inp_block[26-1];
   assign out_block[12] = inp_block[5-1 ];
   assign out_block[13] = inp_block[18-1];   
   assign out_block[14] = inp_block[31-1];
   assign out_block[15] = inp_block[10-1];
   assign out_block[16] = inp_block[2-1 ];
   assign out_block[17] = inp_block[8-1 ];
   assign out_block[18] = inp_block[24-1];
   assign out_block[19] = inp_block[14-1];
   assign out_block[20] = inp_block[32-1];
   assign out_block[21] = inp_block[27-1];
   assign out_block[22] = inp_block[3-1 ];
   assign out_block[23] = inp_block[9-1 ];   
   assign out_block[24] = inp_block[19-1];
   assign out_block[25] = inp_block[13-1];
   assign out_block[26] = inp_block[30-1];
   assign out_block[27] = inp_block[6-1 ];
   assign out_block[28] = inp_block[22-1];
   assign out_block[29] = inp_block[11-1];
   assign out_block[30] = inp_block[4-1 ];
   assign out_block[31] = inp_block[25-1];
 -----/\----- EXCLUDED -----/\----- */
   
endmodule // SF

// Expansion Function
module EF (inp_block, out_block);

   input logic [31:0] inp_block;
   output logic [47:0] out_block;

   assign out_block[ 0] = inp_block[32-1];
   assign out_block[ 1] = inp_block[1-1 ];
   assign out_block[ 2] = inp_block[2-1 ];
   assign out_block[ 3] = inp_block[3-1 ];
   assign out_block[ 4] = inp_block[4-1 ];
   assign out_block[ 5] = inp_block[5-1 ];
   assign out_block[ 6] = inp_block[4-1 ];
   assign out_block[ 7] = inp_block[5-1 ];
   assign out_block[ 8] = inp_block[6-1 ];
   assign out_block[ 9] = inp_block[7-1 ];   
   assign out_block[10] = inp_block[8-1 ];
   assign out_block[11] = inp_block[9-1 ];
   assign out_block[12] = inp_block[8-1 ];
   assign out_block[13] = inp_block[9-1 ];
   assign out_block[14] = inp_block[10-1];
   assign out_block[15] = inp_block[11-1];
   assign out_block[16] = inp_block[12-1];
   assign out_block[17] = inp_block[13-1];
   assign out_block[18] = inp_block[12-1];
   assign out_block[19] = inp_block[13-1];   
   assign out_block[20] = inp_block[14-1];
   assign out_block[21] = inp_block[15-1];
   assign out_block[22] = inp_block[16-1];
   assign out_block[23] = inp_block[17-1];
   assign out_block[24] = inp_block[16-1];
   assign out_block[25] = inp_block[17-1];
   assign out_block[26] = inp_block[18-1];
   assign out_block[27] = inp_block[19-1];
   assign out_block[28] = inp_block[20-1];
   assign out_block[29] = inp_block[21-1];   
   assign out_block[30] = inp_block[20-1];
   assign out_block[31] = inp_block[21-1];
   assign out_block[32] = inp_block[22-1];
   assign out_block[33] = inp_block[23-1];
   assign out_block[34] = inp_block[24-1];
   assign out_block[35] = inp_block[25-1];
   assign out_block[36] = inp_block[24-1];
   assign out_block[37] = inp_block[25-1];
   assign out_block[38] = inp_block[26-1];
   assign out_block[39] = inp_block[27-1];   
   assign out_block[40] = inp_block[28-1];
   assign out_block[41] = inp_block[29-1];
   assign out_block[42] = inp_block[28-1];
   assign out_block[43] = inp_block[29-1];
   assign out_block[44] = inp_block[30-1];
   assign out_block[45] = inp_block[31-1];
   assign out_block[46] = inp_block[32-1];
   assign out_block[47] = inp_block[1-1 ];
   
endmodule // EF

module feistel (inp_block, subkey, out_block);

   input logic [31:0]  inp_block;
   input logic [47:0]  subkey;
   output logic [31:0] out_block;

   logic [47:0]        ep_out;
   logic [47:0]        sbox_pre;   
   logic [3:0] 	       sb1out, sb2out, sb3out, sb4out;
   logic [3:0] 	       sb5out, sb6out, sb7out, sb8out;
   logic [5:0] 	       sb1in, sb2in, sb3in, sb4in;
   logic [5:0] 	       sb5in, sb6in, sb7in, sb8in;      

   // Expansion Function
   EF b1 (inp_block, ep_out);
   // Separate bits for each S-box
   assign sbox_pre = ep_out^subkey;
   assign sb8in = {sbox_pre[5], sbox_pre[0], sbox_pre[4:1]};
   assign sb7in = {sbox_pre[11], sbox_pre[6], sbox_pre[10:7]};
   assign sb6in = {sbox_pre[17], sbox_pre[12], sbox_pre[16:13]};
   assign sb5in = {sbox_pre[23], sbox_pre[18], sbox_pre[22:19]};   
   assign sb4in = {sbox_pre[29], sbox_pre[24], sbox_pre[28:25]};
   assign sb3in = {sbox_pre[35], sbox_pre[30], sbox_pre[34:31]};
   assign sb2in = {sbox_pre[41], sbox_pre[36], sbox_pre[40:37]};
   assign sb1in = {sbox_pre[47], sbox_pre[42], sbox_pre[46:43]};
   // S-boxes
   S1_Box s1 (sb1in, sb1out);
   S2_Box s2 (sb2in, sb2out);
   S3_Box s3 (sb3in, sb3out);
   S4_Box s4 (sb4in, sb4out);   
   S5_Box s5 (sb5in, sb5out);
   S6_Box s6 (sb6in, sb6out);
   S7_Box s7 (sb7in, sb7out);
   S8_Box s8 (sb8in, sb8out);
   // Straight Function
   SF b2 ({sb1out, sb2out, sb3out, sb4out,
	   sb5out, sb6out, sb7out, sb8out},
	  out_block);   
   
endmodule // Feistel

// DES block round
module round (inp_block, subkey, out_block);

   input logic [63:0]  inp_block;
   input logic [47:0]  subkey;
   output logic [63:0] out_block;

   logic [31:0]        Left0;
   logic [31:0]        Right0;
   logic [31:0]        Left1;
   logic [31:0]        Right1;   
   logic [31:0]        f_out;   

   assign {Left0, Right0} = inp_block;
   feistel fk (Right0, subkey, f_out);
   assign Right1 = f_out^Left0;
   assign Left1 = Right0;
   assign out_block = {Left1, Right1};  

endmodule // round1

// Initial Permutation
module IP (inp_block, out_block);

   input logic [63:0]  inp_block;
   output logic [63:0] out_block;

   assign out_block[0] = inp_block[58-1];
   assign out_block[1] = inp_block[50-1];
   assign out_block[2] = inp_block[42-1];
   assign out_block[3] = inp_block[34-1];
   assign out_block[4] = inp_block[26-1];
   assign out_block[5] = inp_block[18-1];
   assign out_block[6] = inp_block[10-1];
   assign out_block[7] = inp_block[2-1 ];
   assign out_block[8] = inp_block[60-1];
   assign out_block[9] = inp_block[52-1];   
   assign out_block[10] = inp_block[44-1];   
   assign out_block[11] = inp_block[36-1];
   assign out_block[12] = inp_block[28-1];
   assign out_block[13] = inp_block[20-1];
   assign out_block[14] = inp_block[12-1];
   assign out_block[15] = inp_block[4-1 ];
   assign out_block[16] = inp_block[62-1];
   assign out_block[17] = inp_block[54-1];
   assign out_block[18] = inp_block[46-1];
   assign out_block[19] = inp_block[38-1];   
   assign out_block[20] = inp_block[30-1];
   assign out_block[21] = inp_block[22-1];   
   assign out_block[22] = inp_block[14-1];
   assign out_block[23] = inp_block[6-1 ];
   assign out_block[24] = inp_block[64-1];
   assign out_block[25] = inp_block[56-1];
   assign out_block[26] = inp_block[48-1];
   assign out_block[27] = inp_block[40-1];
   assign out_block[28] = inp_block[32-1];
   assign out_block[29] = inp_block[24-1];   
   assign out_block[30] = inp_block[16-1];
   assign out_block[31] = inp_block[8-1 ];   
   assign out_block[32] = inp_block[57-1];
   assign out_block[33] = inp_block[49-1];
   assign out_block[34] = inp_block[41-1];
   assign out_block[35] = inp_block[33-1];
   assign out_block[36] = inp_block[25-1];
   assign out_block[37] = inp_block[17-1];
   assign out_block[38] = inp_block[9-1 ];   
   assign out_block[39] = inp_block[1-1 ];   
   assign out_block[40] = inp_block[59-1];
   assign out_block[41] = inp_block[51-1];   
   assign out_block[42] = inp_block[43-1];
   assign out_block[43] = inp_block[35-1];
   assign out_block[44] = inp_block[27-1];
   assign out_block[45] = inp_block[19-1];
   assign out_block[46] = inp_block[11-1];
   assign out_block[47] = inp_block[3-1 ];
   assign out_block[48] = inp_block[61-1];
   assign out_block[49] = inp_block[53-1];   
   assign out_block[50] = inp_block[45-1];
   assign out_block[51] = inp_block[37-1];   
   assign out_block[52] = inp_block[29-1];
   assign out_block[53] = inp_block[21-1];
   assign out_block[54] =  inp_block[13-1];
   assign out_block[55] =  inp_block[5-1 ];
   assign out_block[56] =  inp_block[63-1];
   assign out_block[57] =  inp_block[55-1];
   assign out_block[58] =  inp_block[47-1];
   assign out_block[59] =  inp_block[39-1];   
   assign out_block[60] =  inp_block[31-1];
   assign out_block[61] =  inp_block[23-1];    
   assign out_block[62] =  inp_block[15-1];
   assign out_block[63] =  inp_block[7-1 ];   
   
endmodule // IP

// Final Permutation
module FP (inp_block, out_block);

   input logic [63:0]  inp_block;
   output logic [63:0] out_block;

   assign out_block[ 0] = inp_block[40-1];
   assign out_block[ 1] = inp_block[8-1 ];
   assign out_block[ 2] = inp_block[48-1];
   assign out_block[ 3] = inp_block[16-1];
   assign out_block[ 4] = inp_block[56-1];
   assign out_block[ 5] = inp_block[24-1];
   assign out_block[ 6] = inp_block[64-1];
   assign out_block[ 7] = inp_block[32-1];
   assign out_block[ 8] = inp_block[39-1];
   assign out_block[ 9] = inp_block[7-1 ];   
   assign out_block[10] = inp_block[47-1];   
   assign out_block[11] = inp_block[15-1];
   assign out_block[12] = inp_block[55-1];
   assign out_block[13] = inp_block[23-1];
   assign out_block[14] = inp_block[63-1];
   assign out_block[15] = inp_block[31-1];
   assign out_block[16] = inp_block[38-1];
   assign out_block[17] = inp_block[6-1 ];
   assign out_block[18] = inp_block[46-1];
   assign out_block[19] = inp_block[14-1];   
   assign out_block[20] = inp_block[54-1];
   assign out_block[21] = inp_block[22-1];   
   assign out_block[22] = inp_block[62-1];
   assign out_block[23] = inp_block[30-1];
   assign out_block[24] = inp_block[37-1];
   assign out_block[25] = inp_block[5-1 ];
   assign out_block[26] = inp_block[45-1];
   assign out_block[27] = inp_block[13-1];
   assign out_block[28] = inp_block[53-1];
   assign out_block[29] = inp_block[21-1];   
   assign out_block[30] = inp_block[61-1];
   assign out_block[31] = inp_block[29-1];   
   assign out_block[32] = inp_block[36-1];
   assign out_block[33] = inp_block[4-1 ];
   assign out_block[34] = inp_block[44-1];
   assign out_block[35] = inp_block[12-1];
   assign out_block[36] = inp_block[52-1];
   assign out_block[37] = inp_block[20-1];
   assign out_block[38] = inp_block[60-1];   
   assign out_block[39] = inp_block[28-1];   
   assign out_block[40] = inp_block[35-1];
   assign out_block[41] = inp_block[3-1 ];   
   assign out_block[42] = inp_block[43-1];
   assign out_block[43] = inp_block[11-1];
   assign out_block[44] = inp_block[51-1];
   assign out_block[45] = inp_block[19-1];
   assign out_block[46] = inp_block[59-1];
   assign out_block[47] = inp_block[27-1];
   assign out_block[48] = inp_block[34-1];
   assign out_block[49] = inp_block[2-1 ];   
   assign out_block[50] = inp_block[42-1];
   assign out_block[51] = inp_block[10-1];   
   assign out_block[52] = inp_block[50-1];
   assign out_block[53] = inp_block[18-1];
   assign out_block[54] = inp_block[58-1];
   assign out_block[55] = inp_block[26-1];
   assign out_block[56] = inp_block[33-1];
   assign out_block[57] = inp_block[1-1 ];
   assign out_block[58] = inp_block[41-1];
   assign out_block[59] = inp_block[9-1 ];   
   assign out_block[60] = inp_block[49-1];
   assign out_block[61] = inp_block[17-1];    
   assign out_block[62] = inp_block[57-1];
   assign out_block[63] = inp_block[25-1];   
   
endmodule // round1

module S1_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)             
	  6'd0  : out_bits = 4'd14;             
	  6'd1  : out_bits = 4'd4;             
	  6'd2  : out_bits = 4'd13;            
	  6'd3  : out_bits = 4'd1;             
	  6'd4  : out_bits = 4'd2;             
	  6'd5  : out_bits = 4'd15;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd8;             
	  6'd8  : out_bits = 4'd3;             
	  6'd9  : out_bits = 4'd10;             
	  6'd10 : out_bits = 4'd6;             
	  6'd11 : out_bits = 4'd12;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd9;             
	  6'd14 : out_bits = 4'd0;             
	  6'd15 : out_bits = 4'd7;             
	  6'd16 : out_bits = 4'd0;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd7;             
	  6'd19 : out_bits = 4'd4;             
	  6'd20 : out_bits = 4'd14;             
	  6'd21 : out_bits = 4'd2;             
	  6'd22 : out_bits = 4'd13;             
	  6'd23 : out_bits = 4'd1;             
	  6'd24 : out_bits = 4'd10;             
	  6'd25 : out_bits = 4'd6;             
	  6'd26 : out_bits = 4'd12;             
	  6'd27 : out_bits = 4'd11;             
	  6'd28 : out_bits = 4'd9;             
	  6'd29 : out_bits = 4'd5;             
	  6'd30 : out_bits = 4'd3;             
	  6'd31 : out_bits = 4'd8;             
	  6'd32 : out_bits = 4'd4;             
	  6'd33 : out_bits = 4'd1;             
	  6'd34 : out_bits = 4'd14;             
	  6'd35 : out_bits = 4'd8;             
	  6'd36 : out_bits = 4'd13;             
	  6'd37 : out_bits = 4'd6;             
	  6'd38 : out_bits = 4'd2;             
	  6'd39 : out_bits = 4'd11;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd12;             
	  6'd42 : out_bits = 4'd9;             
	  6'd43 : out_bits = 4'd7;             
	  6'd44 : out_bits = 4'd3;             
	  6'd45 : out_bits = 4'd10;             
	  6'd46 : out_bits = 4'd5;             
	  6'd47 : out_bits = 4'd0;             
	  6'd48 : out_bits = 4'd15;             
	  6'd49 : out_bits = 4'd12;             
	  6'd50 : out_bits = 4'd8;             
	  6'd51 : out_bits = 4'd2;             
	  6'd52 : out_bits = 4'd4;             
	  6'd53 : out_bits = 4'd9;            
	  6'd54 : out_bits = 4'd1;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd5;        
	  6'd57 : out_bits = 4'd11;        
	  6'd58 : out_bits = 4'd3;       
	  6'd59 : out_bits = 4'd14;       
	  6'd60 : out_bits = 4'd10;       
	  6'd61 : out_bits = 4'd0;       
	  6'd62 : out_bits = 4'd6;      
	  6'd63 : out_bits = 4'd13;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S1_Box

module S2_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)             
	  6'd0  : out_bits = 4'd15;             
	  6'd1  : out_bits = 4'd1;             
	  6'd2  : out_bits = 4'd8;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd11;             
	  6'd6  : out_bits = 4'd3;             
	  6'd7  : out_bits = 4'd4;             
	  6'd8  : out_bits = 4'd9;             
	  6'd9  : out_bits = 4'd7;             
	  6'd10 : out_bits = 4'd2;             
	  6'd11 : out_bits = 4'd13;             
	  6'd12 : out_bits = 4'd12;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd5;             
	  6'd15 : out_bits = 4'd10;             
	  6'd16 : out_bits = 4'd3;             
	  6'd17 : out_bits = 4'd13;             
	  6'd18 : out_bits = 4'd4;             
	  6'd19 : out_bits = 4'd7;             
	  6'd20 : out_bits = 4'd15;             
	  6'd21 : out_bits = 4'd2;             
	  6'd22 : out_bits = 4'd8;             
	  6'd23 : out_bits = 4'd14;             
	  6'd24 : out_bits = 4'd12;             
	  6'd25 : out_bits = 4'd0;             
	  6'd26 : out_bits = 4'd1;             
	  6'd27 : out_bits = 4'd10;             
	  6'd28 : out_bits = 4'd6;             
	  6'd29 : out_bits = 4'd9;             
	  6'd30 : out_bits = 4'd11;             
	  6'd31 : out_bits = 4'd5;             
	  6'd32 : out_bits = 4'd0;             
	  6'd33 : out_bits = 4'd14;             
	  6'd34 : out_bits = 4'd7;             
	  6'd35 : out_bits = 4'd11;             
	  6'd36 : out_bits = 4'd10;             
	  6'd37 : out_bits = 4'd4;             
	  6'd38 : out_bits = 4'd13;             
	  6'd39 : out_bits = 4'd1;             
	  6'd40 : out_bits = 4'd5;             
	  6'd41 : out_bits = 4'd8;             
	  6'd42 : out_bits = 4'd12;             
	  6'd43 : out_bits = 4'd6;             
	  6'd44 : out_bits = 4'd9;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd2;             
	  6'd47 : out_bits = 4'd15;             
	  6'd48 : out_bits = 4'd13;             
	  6'd49 : out_bits = 4'd8;             
	  6'd50 : out_bits = 4'd10;             
	  6'd51 : out_bits = 4'd1;             
	  6'd52 : out_bits = 4'd3;             
	  6'd53 : out_bits = 4'd15;            
	  6'd54 : out_bits = 4'd4;             
	  6'd55 : out_bits = 4'd2;            
	  6'd56 : out_bits = 4'd11;        
	  6'd57 : out_bits = 4'd6;        
	  6'd58 : out_bits = 4'd7;       
	  6'd59 : out_bits = 4'd12;       
	  6'd60 : out_bits = 4'd0;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd14;      
	  6'd63 : out_bits = 4'd9;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S2_Box

module S3_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)
	  6'd0  : out_bits = 4'd10;             
	  6'd1  : out_bits = 4'd0;             
	  6'd2  : out_bits = 4'd9;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd3;             
	  6'd6  : out_bits = 4'd15;             
	  6'd7  : out_bits = 4'd5;             
	  6'd8  : out_bits = 4'd1;             
	  6'd9  : out_bits = 4'd13;             
	  6'd10 : out_bits = 4'd12;             
	  6'd11 : out_bits = 4'd7;             
	  6'd12 : out_bits = 4'd11;             
	  6'd13 : out_bits = 4'd4;             
	  6'd14 : out_bits = 4'd2;             
	  6'd15 : out_bits = 4'd8;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd7;             
	  6'd18 : out_bits = 4'd0;             
	  6'd19 : out_bits = 4'd9;             
	  6'd20 : out_bits = 4'd3;             
	  6'd21 : out_bits = 4'd4;             
	  6'd22 : out_bits = 4'd6;             
	  6'd23 : out_bits = 4'd10;             
	  6'd24 : out_bits = 4'd2;             
	  6'd25 : out_bits = 4'd8;             
	  6'd26 : out_bits = 4'd5;             
	  6'd27 : out_bits = 4'd14;             
	  6'd28 : out_bits = 4'd12;             
	  6'd29 : out_bits = 4'd11;             
	  6'd30 : out_bits = 4'd15;             
	  6'd31 : out_bits = 4'd1;             
	  6'd32 : out_bits = 4'd13;             
	  6'd33 : out_bits = 4'd6;             
	  6'd34 : out_bits = 4'd4;             
	  6'd35 : out_bits = 4'd9;             
	  6'd36 : out_bits = 4'd8;             
	  6'd37 : out_bits = 4'd15;             
	  6'd38 : out_bits = 4'd3;             
	  6'd39 : out_bits = 4'd0;             
	  6'd40 : out_bits = 4'd11;             
	  6'd41 : out_bits = 4'd1;             
	  6'd42 : out_bits = 4'd2;             
	  6'd43 : out_bits = 4'd12;             
	  6'd44 : out_bits = 4'd5;             
	  6'd45 : out_bits = 4'd10;             
	  6'd46 : out_bits = 4'd14;             
	  6'd47 : out_bits = 4'd7;             
	  6'd48 : out_bits = 4'd1;             
	  6'd49 : out_bits = 4'd10;             
	  6'd50 : out_bits = 4'd13;             
	  6'd51 : out_bits = 4'd0;             
	  6'd52 : out_bits = 4'd6;             
	  6'd53 : out_bits = 4'd9;            
	  6'd54 : out_bits = 4'd8;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd4;        
	  6'd57 : out_bits = 4'd15;        
	  6'd58 : out_bits = 4'd14;       
	  6'd59 : out_bits = 4'd3;       
	  6'd60 : out_bits = 4'd11;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd2;      
	  6'd63 : out_bits = 4'd12;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S3_Box

module S4_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)   
	  6'd0  : out_bits = 4'd7;             
	  6'd1  : out_bits = 4'd13;             
	  6'd2  : out_bits = 4'd14;            
	  6'd3  : out_bits = 4'd3;             
	  6'd4  : out_bits = 4'd0;             
	  6'd5  : out_bits = 4'd6;             
	  6'd6  : out_bits = 4'd9;             
	  6'd7  : out_bits = 4'd10;             
	  6'd8  : out_bits = 4'd1;             
	  6'd9  : out_bits = 4'd2;             
	  6'd10 : out_bits = 4'd8;             
	  6'd11 : out_bits = 4'd5;             
	  6'd12 : out_bits = 4'd11;             
	  6'd13 : out_bits = 4'd12;             
	  6'd14 : out_bits = 4'd4;             
	  6'd15 : out_bits = 4'd15;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd8;             
	  6'd18 : out_bits = 4'd11;             
	  6'd19 : out_bits = 4'd5;             
	  6'd20 : out_bits = 4'd6;             
	  6'd21 : out_bits = 4'd15;             
	  6'd22 : out_bits = 4'd0;             
	  6'd23 : out_bits = 4'd3;             
	  6'd24 : out_bits = 4'd4;             
	  6'd25 : out_bits = 4'd7;             
	  6'd26 : out_bits = 4'd2;             
	  6'd27 : out_bits = 4'd12;             
	  6'd28 : out_bits = 4'd1;             
	  6'd29 : out_bits = 4'd10;             
	  6'd30 : out_bits = 4'd14;             
	  6'd31 : out_bits = 4'd9;             
	  6'd32 : out_bits = 4'd10;             
	  6'd33 : out_bits = 4'd6;             
	  6'd34 : out_bits = 4'd9;             
	  6'd35 : out_bits = 4'd0;             
	  6'd36 : out_bits = 4'd12;             
	  6'd37 : out_bits = 4'd11;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd13;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd1;             
	  6'd42 : out_bits = 4'd3;             
	  6'd43 : out_bits = 4'd14;             
	  6'd44 : out_bits = 4'd5;             
	  6'd45 : out_bits = 4'd2;             
	  6'd46 : out_bits = 4'd8;             
	  6'd47 : out_bits = 4'd4;             
	  6'd48 : out_bits = 4'd3;             
	  6'd49 : out_bits = 4'd15;             
	  6'd50 : out_bits = 4'd0;             
	  6'd51 : out_bits = 4'd6;             
	  6'd52 : out_bits = 4'd10;             
	  6'd53 : out_bits = 4'd1;            
	  6'd54 : out_bits = 4'd13;             
	  6'd55 : out_bits = 4'd8;            
	  6'd56 : out_bits = 4'd9;        
	  6'd57 : out_bits = 4'd4;        
	  6'd58 : out_bits = 4'd5;       
	  6'd59 : out_bits = 4'd11;       
	  6'd60 : out_bits = 4'd12;       
	  6'd61 : out_bits = 4'd7;       
	  6'd62 : out_bits = 4'd2;      
	  6'd63 : out_bits = 4'd14;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S4_Box

module S5_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)   
	  6'd0  : out_bits = 4'd2;             
	  6'd1  : out_bits = 4'd12;             
	  6'd2  : out_bits = 4'd4;            
	  6'd3  : out_bits = 4'd1;             
	  6'd4  : out_bits = 4'd7;             
	  6'd5  : out_bits = 4'd10;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd6;             
	  6'd8  : out_bits = 4'd8;             
	  6'd9  : out_bits = 4'd5;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd15;             
	  6'd12 : out_bits = 4'd13;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd14;             
	  6'd15 : out_bits = 4'd9;             
	  6'd16 : out_bits = 4'd14;             
	  6'd17 : out_bits = 4'd11;             
	  6'd18 : out_bits = 4'd2;             
	  6'd19 : out_bits = 4'd12;             
	  6'd20 : out_bits = 4'd4;             
	  6'd21 : out_bits = 4'd7;             
	  6'd22 : out_bits = 4'd13;             
	  6'd23 : out_bits = 4'd1;             
	  6'd24 : out_bits = 4'd5;             
	  6'd25 : out_bits = 4'd0;             
	  6'd26 : out_bits = 4'd15;             
	  6'd27 : out_bits = 4'd10;             
	  6'd28 : out_bits = 4'd3;             
	  6'd29 : out_bits = 4'd9;             
	  6'd30 : out_bits = 4'd8;             
	  6'd31 : out_bits = 4'd6;             
	  6'd32 : out_bits = 4'd4;             
	  6'd33 : out_bits = 4'd2;             
	  6'd34 : out_bits = 4'd1;             
	  6'd35 : out_bits = 4'd11;             
	  6'd36 : out_bits = 4'd10;             
	  6'd37 : out_bits = 4'd13;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd8;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd9;             
	  6'd42 : out_bits = 4'd12;             
	  6'd43 : out_bits = 4'd5;             
	  6'd44 : out_bits = 4'd6;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd0;             
	  6'd47 : out_bits = 4'd14;             
	  6'd48 : out_bits = 4'd11;             
	  6'd49 : out_bits = 4'd8;             
	  6'd50 : out_bits = 4'd12;             
	  6'd51 : out_bits = 4'd7;             
	  6'd52 : out_bits = 4'd1;             
	  6'd53 : out_bits = 4'd14;            
	  6'd54 : out_bits = 4'd2;             
	  6'd55 : out_bits = 4'd13;            
	  6'd56 : out_bits = 4'd6;        
	  6'd57 : out_bits = 4'd15;        
	  6'd58 : out_bits = 4'd0;       
	  6'd59 : out_bits = 4'd9;       
	  6'd60 : out_bits = 4'd10;       
	  6'd61 : out_bits = 4'd4;       
	  6'd62 : out_bits = 4'd5;      
	  6'd63 : out_bits = 4'd3;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S5_Box

module S6_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)   
	  6'd0  : out_bits = 4'd12;             
	  6'd1  : out_bits = 4'd1;             
	  6'd2  : out_bits = 4'd10;            
	  6'd3  : out_bits = 4'd15;             
	  6'd4  : out_bits = 4'd9;             
	  6'd5  : out_bits = 4'd2;             
	  6'd6  : out_bits = 4'd6;             
	  6'd7  : out_bits = 4'd8;             
	  6'd8  : out_bits = 4'd0;             
	  6'd9  : out_bits = 4'd13;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd4;             
	  6'd12 : out_bits = 4'd14;             
	  6'd13 : out_bits = 4'd7;             
	  6'd14 : out_bits = 4'd5;             
	  6'd15 : out_bits = 4'd11;             
	  6'd16 : out_bits = 4'd10;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd4;             
	  6'd19 : out_bits = 4'd2;             
	  6'd20 : out_bits = 4'd7;             
	  6'd21 : out_bits = 4'd12;             
	  6'd22 : out_bits = 4'd9;             
	  6'd23 : out_bits = 4'd5;             
	  6'd24 : out_bits = 4'd6;             
	  6'd25 : out_bits = 4'd1;             
	  6'd26 : out_bits = 4'd13;             
	  6'd27 : out_bits = 4'd14;             
	  6'd28 : out_bits = 4'd0;             
	  6'd29 : out_bits = 4'd11;             
	  6'd30 : out_bits = 4'd3;             
	  6'd31 : out_bits = 4'd8;             
	  6'd32 : out_bits = 4'd9;             
	  6'd33 : out_bits = 4'd14;             
	  6'd34 : out_bits = 4'd15;             
	  6'd35 : out_bits = 4'd5;             
	  6'd36 : out_bits = 4'd2;             
	  6'd37 : out_bits = 4'd8;             
	  6'd38 : out_bits = 4'd12;             
	  6'd39 : out_bits = 4'd3;             
	  6'd40 : out_bits = 4'd7;             
	  6'd41 : out_bits = 4'd0;             
	  6'd42 : out_bits = 4'd4;             
	  6'd43 : out_bits = 4'd10;             
	  6'd44 : out_bits = 4'd1;             
	  6'd45 : out_bits = 4'd13;             
	  6'd46 : out_bits = 4'd11;             
	  6'd47 : out_bits = 4'd6;             
	  6'd48 : out_bits = 4'd4;             
	  6'd49 : out_bits = 4'd3;             
	  6'd50 : out_bits = 4'd2;             
	  6'd51 : out_bits = 4'd12;             
	  6'd52 : out_bits = 4'd9;             
	  6'd53 : out_bits = 4'd5;            
	  6'd54 : out_bits = 4'd15;             
	  6'd55 : out_bits = 4'd10;            
	  6'd56 : out_bits = 4'd11;        
	  6'd57 : out_bits = 4'd14;        
	  6'd58 : out_bits = 4'd1;       
	  6'd59 : out_bits = 4'd7;       
	  6'd60 : out_bits = 4'd6;       
	  6'd61 : out_bits = 4'd0;       
	  6'd62 : out_bits = 4'd8;      
	  6'd63 : out_bits = 4'd13;	  
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S6_Box

module S7_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)   
	  6'd0  : out_bits = 4'd4;             
	  6'd1  : out_bits = 4'd11;             
	  6'd2  : out_bits = 4'd2;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd15;             
	  6'd5  : out_bits = 4'd0;             
	  6'd6  : out_bits = 4'd8;             
	  6'd7  : out_bits = 4'd13;             
	  6'd8  : out_bits = 4'd3;             
	  6'd9  : out_bits = 4'd12;             
	  6'd10 : out_bits = 4'd9;             
	  6'd11 : out_bits = 4'd7;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd10;             
	  6'd14 : out_bits = 4'd6;             
	  6'd15 : out_bits = 4'd1;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd0;             
	  6'd18 : out_bits = 4'd11;             
	  6'd19 : out_bits = 4'd7;             
	  6'd20 : out_bits = 4'd4;             
	  6'd21 : out_bits = 4'd9;             
	  6'd22 : out_bits = 4'd1;             
	  6'd23 : out_bits = 4'd10;             
	  6'd24 : out_bits = 4'd14;             
	  6'd25 : out_bits = 4'd3;             
	  6'd26 : out_bits = 4'd5;             
	  6'd27 : out_bits = 4'd12;             
	  6'd28 : out_bits = 4'd2;             
	  6'd29 : out_bits = 4'd15;             
	  6'd30 : out_bits = 4'd8;             
	  6'd31 : out_bits = 4'd6;             
	  6'd32 : out_bits = 4'd1;             
	  6'd33 : out_bits = 4'd4;             
	  6'd34 : out_bits = 4'd11;             
	  6'd35 : out_bits = 4'd13;             
	  6'd36 : out_bits = 4'd12;             
	  6'd37 : out_bits = 4'd3;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd14;             
	  6'd40 : out_bits = 4'd10;             
	  6'd41 : out_bits = 4'd15;             
	  6'd42 : out_bits = 4'd6;             
	  6'd43 : out_bits = 4'd8;             
	  6'd44 : out_bits = 4'd0;             
	  6'd45 : out_bits = 4'd5;             
	  6'd46 : out_bits = 4'd9;             
	  6'd47 : out_bits = 4'd2;             
	  6'd48 : out_bits = 4'd6;             
	  6'd49 : out_bits = 4'd11;             
	  6'd50 : out_bits = 4'd13;             
	  6'd51 : out_bits = 4'd8;             
	  6'd52 : out_bits = 4'd1;             
	  6'd53 : out_bits = 4'd4;            
	  6'd54 : out_bits = 4'd10;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd9;        
	  6'd57 : out_bits = 4'd5;        
	  6'd58 : out_bits = 4'd0;       
	  6'd59 : out_bits = 4'd15;       
	  6'd60 : out_bits = 4'd14;       
	  6'd61 : out_bits = 4'd2;       
	  6'd62 : out_bits = 4'd3;      
	  6'd63 : out_bits = 4'd12;  
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S7_Box

module S8_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case (inp_bits)   
	  6'd0  : out_bits = 4'd13;             
	  6'd1  : out_bits = 4'd2;             
	  6'd2  : out_bits = 4'd8;            
	  6'd3  : out_bits = 4'd4;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd15;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd1;             
	  6'd8  : out_bits = 4'd10;             
	  6'd9  : out_bits = 4'd9;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd14;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd12;             
	  6'd15 : out_bits = 4'd7;             
	  6'd16 : out_bits = 4'd1;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd13;             
	  6'd19 : out_bits = 4'd8;             
	  6'd20 : out_bits = 4'd10;             
	  6'd21 : out_bits = 4'd3;             
	  6'd22 : out_bits = 4'd7;             
	  6'd23 : out_bits = 4'd4;             
	  6'd24 : out_bits = 4'd12;             
	  6'd25 : out_bits = 4'd5;             
	  6'd26 : out_bits = 4'd6;             
	  6'd27 : out_bits = 4'd11;             
	  6'd28 : out_bits = 4'd0;             
	  6'd29 : out_bits = 4'd14;             
	  6'd30 : out_bits = 4'd9;             
	  6'd31 : out_bits = 4'd2;             
	  6'd32 : out_bits = 4'd7;             
	  6'd33 : out_bits = 4'd11;             
	  6'd34 : out_bits = 4'd4;             
	  6'd35 : out_bits = 4'd1;             
	  6'd36 : out_bits = 4'd9;             
	  6'd37 : out_bits = 4'd12;             
	  6'd38 : out_bits = 4'd14;             
	  6'd39 : out_bits = 4'd2;             
	  6'd40 : out_bits = 4'd0;             
	  6'd41 : out_bits = 4'd6;             
	  6'd42 : out_bits = 4'd10;             
	  6'd43 : out_bits = 4'd13;             
	  6'd44 : out_bits = 4'd15;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd5;             
	  6'd47 : out_bits = 4'd8;             
	  6'd48 : out_bits = 4'd2;             
	  6'd49 : out_bits = 4'd1;             
	  6'd50 : out_bits = 4'd14;             
	  6'd51 : out_bits = 4'd7;             
	  6'd52 : out_bits = 4'd4;             
	  6'd53 : out_bits = 4'd10;            
	  6'd54 : out_bits = 4'd8;             
	  6'd55 : out_bits = 4'd13;            
	  6'd56 : out_bits = 4'd15;        
	  6'd57 : out_bits = 4'd12;        
	  6'd58 : out_bits = 4'd9;       
	  6'd59 : out_bits = 4'd0;       
	  6'd60 : out_bits = 4'd3;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd6;      
	  6'd63 : out_bits = 4'd11;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S8_Box

module DES (input logic [63:0] key, input logic [63:0] plaintext, 
	    input logic encrypt, output logic [63:0] ciphertext);

   logic [47:0] 	SubKey1, SubKey2, SubKey3, SubKey4;   
   logic [47:0] 	SubKey5, SubKey6, SubKey7, SubKey8;   
   logic [47:0] 	SubKey9, SubKey10, SubKey11, SubKey12;
   logic [47:0] 	SubKey13, SubKey14, SubKey15, SubKey16;
   logic [63:0] 	ip_out;
   logic [63:0] 	r1_out, r2_out, r3_out, r4_out;
   logic [63:0] 	r5_out, r6_out, r7_out, r8_out;
   logic [63:0] 	r9_out, r10_out, r11_out, r12_out;
   logic [63:0] 	r13_out, r14_out, r15_out, r16_out;      

   // SubKey generation
   GenerateKeys k1 (key, SubKey1, SubKey2, SubKey3, SubKey4,
		    SubKey5, SubKey6, SubKey7, SubKey8,
		    SubKey9, SubKey10, SubKey11, SubKey12,
		    SubKey13, SubKey14, SubKey15, SubKey16);

   // DES Function
   
   // Initial Permutation
   IP b1 (plaintext, ip_out);
   // round 1
   round b2 (ip_out, SubKey1, r1_out);
   // round 2
   round b3 (r1_out, SubKey2, r2_out);
   // round 3
   round b4 (r2_out, SubKey3, r3_out);
   // round 4
   round b5 (r3_out, SubKey4, r4_out);
   // round 5
   round b6 (r4_out, SubKey5, r5_out);
   // round 6
   round b7 (r5_out, SubKey6, r6_out);
   // round 7
   round b8 (r6_out, SubKey7, r7_out);
   // round 8
   round b9 (r7_out, SubKey8, r8_out);
   // round 9
   round b10 (r8_out, SubKey9, r9_out);
   // round 10
   round b11 (r9_out, SubKey10, r10_out);
   // round 11
   round b12 (r10_out, SubKey11, r11_out);
   // round 12
   round b13 (r11_out, SubKey12, r12_out);
   // round 13
   round b14 (r12_out, SubKey13, r13_out);
   // round 14
   round b15 (r13_out, SubKey14, r14_out);
   // round 15
   round b16 (r14_out, SubKey15, r15_out);
   // round 16
   round b17 (r15_out, SubKey16, r16_out);

   FP FP({r16_out[31:0], r16_out[63:32]}, ciphertext);
  
  // assign ciphertext = r16_out;   
   
endmodule // DES


